magic
tech sky130A
timestamp 1654928256
<< metal3 >>
rect -408 16 408 30
rect -408 -16 -396 16
rect -364 -16 -356 16
rect -324 -16 -316 16
rect -284 -16 -276 16
rect -244 -16 -236 16
rect -204 -16 -196 16
rect -164 -16 -156 16
rect -124 -16 -116 16
rect -84 -16 -76 16
rect -44 -16 -36 16
rect -4 -16 4 16
rect 36 -16 44 16
rect 76 -16 84 16
rect 116 -16 124 16
rect 156 -16 164 16
rect 196 -16 204 16
rect 236 -16 244 16
rect 276 -16 284 16
rect 316 -16 324 16
rect 356 -16 364 16
rect 396 -16 408 16
rect -408 -30 408 -16
<< via3 >>
rect -396 -16 -364 16
rect -356 -16 -324 16
rect -316 -16 -284 16
rect -276 -16 -244 16
rect -236 -16 -204 16
rect -196 -16 -164 16
rect -156 -16 -124 16
rect -116 -16 -84 16
rect -76 -16 -44 16
rect -36 -16 -4 16
rect 4 -16 36 16
rect 44 -16 76 16
rect 84 -16 116 16
rect 124 -16 156 16
rect 164 -16 196 16
rect 204 -16 236 16
rect 244 -16 276 16
rect 284 -16 316 16
rect 324 -16 356 16
rect 364 -16 396 16
<< metal4 >>
rect -408 16 408 30
rect -408 -16 -396 16
rect -364 -16 -356 16
rect -324 -16 -316 16
rect -284 -16 -276 16
rect -244 -16 -236 16
rect -204 -16 -196 16
rect -164 -16 -156 16
rect -124 -16 -116 16
rect -84 -16 -76 16
rect -44 -16 -36 16
rect -4 -16 4 16
rect 36 -16 44 16
rect 76 -16 84 16
rect 116 -16 124 16
rect 156 -16 164 16
rect 196 -16 204 16
rect 236 -16 244 16
rect 276 -16 284 16
rect 316 -16 324 16
rect 356 -16 364 16
rect 396 -16 408 16
rect -408 -30 408 -16
<< end >>
