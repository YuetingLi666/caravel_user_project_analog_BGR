magic
tech sky130A
magscale 1 2
timestamp 1654928256
<< pwell >>
rect 1026 764 1694 996
<< psubdiff >>
rect 1052 931 1668 970
rect 1052 829 1139 931
rect 1581 829 1668 931
rect 1052 790 1668 829
<< psubdiffcont >>
rect 1139 829 1581 931
<< xpolycontact >>
rect 140 1075 572 1645
rect 2148 1075 2580 1645
rect 140 115 572 685
rect 2148 115 2580 685
<< xpolyres >>
rect 572 1075 2148 1645
rect 572 115 2148 685
<< locali >>
rect 140 1897 2580 1910
rect 140 1863 323 1897
rect 357 1863 523 1897
rect 557 1863 723 1897
rect 757 1863 923 1897
rect 957 1863 1123 1897
rect 1157 1863 1323 1897
rect 1357 1863 1523 1897
rect 1557 1863 1723 1897
rect 1757 1863 1923 1897
rect 1957 1863 2123 1897
rect 2157 1863 2323 1897
rect 2357 1863 2580 1897
rect 140 1850 2580 1863
rect 1052 931 1668 970
rect 1052 829 1139 931
rect 1581 829 1668 931
rect 1052 30 1668 829
rect 2148 685 2580 1075
rect 140 17 2580 30
rect 140 -17 323 17
rect 357 -17 523 17
rect 557 -17 723 17
rect 757 -17 923 17
rect 957 -17 1123 17
rect 1157 -17 1323 17
rect 1357 -17 1523 17
rect 1557 -17 1723 17
rect 1757 -17 1923 17
rect 1957 -17 2123 17
rect 2157 -17 2323 17
rect 2357 -17 2580 17
rect 140 -30 2580 -17
<< viali >>
rect 323 1863 357 1897
rect 523 1863 557 1897
rect 723 1863 757 1897
rect 923 1863 957 1897
rect 1123 1863 1157 1897
rect 1323 1863 1357 1897
rect 1523 1863 1557 1897
rect 1723 1863 1757 1897
rect 1923 1863 1957 1897
rect 2123 1863 2157 1897
rect 2323 1863 2357 1897
rect 159 1091 553 1629
rect 2166 1091 2560 1629
rect 159 131 553 669
rect 2166 131 2560 669
rect 323 -17 357 17
rect 523 -17 557 17
rect 723 -17 757 17
rect 923 -17 957 17
rect 1123 -17 1157 17
rect 1323 -17 1357 17
rect 1523 -17 1557 17
rect 1723 -17 1757 17
rect 1923 -17 1957 17
rect 2123 -17 2157 17
rect 2323 -17 2357 17
<< metal1 >>
rect 140 1897 2580 1940
rect 140 1863 323 1897
rect 357 1863 523 1897
rect 557 1863 723 1897
rect 757 1863 923 1897
rect 957 1863 1123 1897
rect 1157 1863 1323 1897
rect 1357 1863 1523 1897
rect 1557 1863 1723 1897
rect 1757 1863 1923 1897
rect 1957 1863 2123 1897
rect 2157 1863 2323 1897
rect 2357 1863 2580 1897
rect 140 1820 2580 1863
rect 151 1629 561 1641
rect 151 1091 159 1629
rect 553 1091 561 1629
rect 151 1079 561 1091
rect 2159 1629 2569 1641
rect 2159 1091 2166 1629
rect 2560 1091 2569 1629
rect 2159 1079 2569 1091
rect 151 669 561 681
rect 151 131 159 669
rect 553 131 561 669
rect 151 119 561 131
rect 2148 669 2580 1079
rect 2148 131 2166 669
rect 2560 131 2580 669
rect 2148 115 2580 131
rect 140 17 2580 60
rect 140 -17 323 17
rect 357 -17 523 17
rect 557 -17 723 17
rect 757 -17 923 17
rect 957 -17 1123 17
rect 1157 -17 1323 17
rect 1357 -17 1523 17
rect 1557 -17 1723 17
rect 1757 -17 1923 17
rect 1957 -17 2123 17
rect 2157 -17 2323 17
rect 2357 -17 2580 17
rect 140 -60 2580 -17
<< labels >>
flabel metal1 s 260 1300 380 1420 1 FreeSans 750 0 0 0 Rin
port 1 nsew
flabel metal1 s 260 340 380 460 1 FreeSans 750 0 0 0 Rout
port 2 nsew
flabel metal1 s 140 1850 200 1910 1 FreeSans 1250 0 0 0 VPWR
port 3 nsew
flabel metal1 s 140 -30 200 30 1 FreeSans 1250 0 0 0 VGND
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2720 1880
<< end >>
