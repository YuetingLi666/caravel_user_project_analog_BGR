magic
tech sky130A
magscale 1 2
timestamp 1655816534
<< nwell >>
rect 120 1707 5842 1940
rect 120 294 5843 1707
rect 217 293 5843 294
<< pmoslvt >>
rect 311 355 711 1645
rect 769 355 1169 1645
rect 1227 355 1627 1645
rect 1685 355 2085 1645
rect 2143 355 2543 1645
rect 2601 355 3001 1645
rect 3059 355 3459 1645
rect 3517 355 3917 1645
rect 3975 355 4375 1645
rect 4433 355 4833 1645
rect 4891 355 5291 1645
rect 5349 355 5749 1645
<< pdiff >>
rect 253 1629 311 1645
rect 253 1595 265 1629
rect 299 1595 311 1629
rect 253 1561 311 1595
rect 253 1527 265 1561
rect 299 1527 311 1561
rect 253 1493 311 1527
rect 253 1459 265 1493
rect 299 1459 311 1493
rect 253 1425 311 1459
rect 253 1391 265 1425
rect 299 1391 311 1425
rect 253 1357 311 1391
rect 253 1323 265 1357
rect 299 1323 311 1357
rect 253 1289 311 1323
rect 253 1255 265 1289
rect 299 1255 311 1289
rect 253 1221 311 1255
rect 253 1187 265 1221
rect 299 1187 311 1221
rect 253 1153 311 1187
rect 253 1119 265 1153
rect 299 1119 311 1153
rect 253 1085 311 1119
rect 253 1051 265 1085
rect 299 1051 311 1085
rect 253 1017 311 1051
rect 253 983 265 1017
rect 299 983 311 1017
rect 253 949 311 983
rect 253 915 265 949
rect 299 915 311 949
rect 253 881 311 915
rect 253 847 265 881
rect 299 847 311 881
rect 253 813 311 847
rect 253 779 265 813
rect 299 779 311 813
rect 253 745 311 779
rect 253 711 265 745
rect 299 711 311 745
rect 253 677 311 711
rect 253 643 265 677
rect 299 643 311 677
rect 253 609 311 643
rect 253 575 265 609
rect 299 575 311 609
rect 253 541 311 575
rect 253 507 265 541
rect 299 507 311 541
rect 253 473 311 507
rect 253 439 265 473
rect 299 439 311 473
rect 253 405 311 439
rect 253 371 265 405
rect 299 371 311 405
rect 253 355 311 371
rect 711 1629 769 1645
rect 711 1595 723 1629
rect 757 1595 769 1629
rect 711 1561 769 1595
rect 711 1527 723 1561
rect 757 1527 769 1561
rect 711 1493 769 1527
rect 711 1459 723 1493
rect 757 1459 769 1493
rect 711 1425 769 1459
rect 711 1391 723 1425
rect 757 1391 769 1425
rect 711 1357 769 1391
rect 711 1323 723 1357
rect 757 1323 769 1357
rect 711 1289 769 1323
rect 711 1255 723 1289
rect 757 1255 769 1289
rect 711 1221 769 1255
rect 711 1187 723 1221
rect 757 1187 769 1221
rect 711 1153 769 1187
rect 711 1119 723 1153
rect 757 1119 769 1153
rect 711 1085 769 1119
rect 711 1051 723 1085
rect 757 1051 769 1085
rect 711 1017 769 1051
rect 711 983 723 1017
rect 757 983 769 1017
rect 711 949 769 983
rect 711 915 723 949
rect 757 915 769 949
rect 711 881 769 915
rect 711 847 723 881
rect 757 847 769 881
rect 711 813 769 847
rect 711 779 723 813
rect 757 779 769 813
rect 711 745 769 779
rect 711 711 723 745
rect 757 711 769 745
rect 711 677 769 711
rect 711 643 723 677
rect 757 643 769 677
rect 711 609 769 643
rect 711 575 723 609
rect 757 575 769 609
rect 711 541 769 575
rect 711 507 723 541
rect 757 507 769 541
rect 711 473 769 507
rect 711 439 723 473
rect 757 439 769 473
rect 711 405 769 439
rect 711 371 723 405
rect 757 371 769 405
rect 711 355 769 371
rect 1169 1629 1227 1645
rect 1169 1595 1181 1629
rect 1215 1595 1227 1629
rect 1169 1561 1227 1595
rect 1169 1527 1181 1561
rect 1215 1527 1227 1561
rect 1169 1493 1227 1527
rect 1169 1459 1181 1493
rect 1215 1459 1227 1493
rect 1169 1425 1227 1459
rect 1169 1391 1181 1425
rect 1215 1391 1227 1425
rect 1169 1357 1227 1391
rect 1169 1323 1181 1357
rect 1215 1323 1227 1357
rect 1169 1289 1227 1323
rect 1169 1255 1181 1289
rect 1215 1255 1227 1289
rect 1169 1221 1227 1255
rect 1169 1187 1181 1221
rect 1215 1187 1227 1221
rect 1169 1153 1227 1187
rect 1169 1119 1181 1153
rect 1215 1119 1227 1153
rect 1169 1085 1227 1119
rect 1169 1051 1181 1085
rect 1215 1051 1227 1085
rect 1169 1017 1227 1051
rect 1169 983 1181 1017
rect 1215 983 1227 1017
rect 1169 949 1227 983
rect 1169 915 1181 949
rect 1215 915 1227 949
rect 1169 881 1227 915
rect 1169 847 1181 881
rect 1215 847 1227 881
rect 1169 813 1227 847
rect 1169 779 1181 813
rect 1215 779 1227 813
rect 1169 745 1227 779
rect 1169 711 1181 745
rect 1215 711 1227 745
rect 1169 677 1227 711
rect 1169 643 1181 677
rect 1215 643 1227 677
rect 1169 609 1227 643
rect 1169 575 1181 609
rect 1215 575 1227 609
rect 1169 541 1227 575
rect 1169 507 1181 541
rect 1215 507 1227 541
rect 1169 473 1227 507
rect 1169 439 1181 473
rect 1215 439 1227 473
rect 1169 405 1227 439
rect 1169 371 1181 405
rect 1215 371 1227 405
rect 1169 355 1227 371
rect 1627 1629 1685 1645
rect 1627 1595 1639 1629
rect 1673 1595 1685 1629
rect 1627 1561 1685 1595
rect 1627 1527 1639 1561
rect 1673 1527 1685 1561
rect 1627 1493 1685 1527
rect 1627 1459 1639 1493
rect 1673 1459 1685 1493
rect 1627 1425 1685 1459
rect 1627 1391 1639 1425
rect 1673 1391 1685 1425
rect 1627 1357 1685 1391
rect 1627 1323 1639 1357
rect 1673 1323 1685 1357
rect 1627 1289 1685 1323
rect 1627 1255 1639 1289
rect 1673 1255 1685 1289
rect 1627 1221 1685 1255
rect 1627 1187 1639 1221
rect 1673 1187 1685 1221
rect 1627 1153 1685 1187
rect 1627 1119 1639 1153
rect 1673 1119 1685 1153
rect 1627 1085 1685 1119
rect 1627 1051 1639 1085
rect 1673 1051 1685 1085
rect 1627 1017 1685 1051
rect 1627 983 1639 1017
rect 1673 983 1685 1017
rect 1627 949 1685 983
rect 1627 915 1639 949
rect 1673 915 1685 949
rect 1627 881 1685 915
rect 1627 847 1639 881
rect 1673 847 1685 881
rect 1627 813 1685 847
rect 1627 779 1639 813
rect 1673 779 1685 813
rect 1627 745 1685 779
rect 1627 711 1639 745
rect 1673 711 1685 745
rect 1627 677 1685 711
rect 1627 643 1639 677
rect 1673 643 1685 677
rect 1627 609 1685 643
rect 1627 575 1639 609
rect 1673 575 1685 609
rect 1627 541 1685 575
rect 1627 507 1639 541
rect 1673 507 1685 541
rect 1627 473 1685 507
rect 1627 439 1639 473
rect 1673 439 1685 473
rect 1627 405 1685 439
rect 1627 371 1639 405
rect 1673 371 1685 405
rect 1627 355 1685 371
rect 2085 1629 2143 1645
rect 2085 1595 2097 1629
rect 2131 1595 2143 1629
rect 2085 1561 2143 1595
rect 2085 1527 2097 1561
rect 2131 1527 2143 1561
rect 2085 1493 2143 1527
rect 2085 1459 2097 1493
rect 2131 1459 2143 1493
rect 2085 1425 2143 1459
rect 2085 1391 2097 1425
rect 2131 1391 2143 1425
rect 2085 1357 2143 1391
rect 2085 1323 2097 1357
rect 2131 1323 2143 1357
rect 2085 1289 2143 1323
rect 2085 1255 2097 1289
rect 2131 1255 2143 1289
rect 2085 1221 2143 1255
rect 2085 1187 2097 1221
rect 2131 1187 2143 1221
rect 2085 1153 2143 1187
rect 2085 1119 2097 1153
rect 2131 1119 2143 1153
rect 2085 1085 2143 1119
rect 2085 1051 2097 1085
rect 2131 1051 2143 1085
rect 2085 1017 2143 1051
rect 2085 983 2097 1017
rect 2131 983 2143 1017
rect 2085 949 2143 983
rect 2085 915 2097 949
rect 2131 915 2143 949
rect 2085 881 2143 915
rect 2085 847 2097 881
rect 2131 847 2143 881
rect 2085 813 2143 847
rect 2085 779 2097 813
rect 2131 779 2143 813
rect 2085 745 2143 779
rect 2085 711 2097 745
rect 2131 711 2143 745
rect 2085 677 2143 711
rect 2085 643 2097 677
rect 2131 643 2143 677
rect 2085 609 2143 643
rect 2085 575 2097 609
rect 2131 575 2143 609
rect 2085 541 2143 575
rect 2085 507 2097 541
rect 2131 507 2143 541
rect 2085 473 2143 507
rect 2085 439 2097 473
rect 2131 439 2143 473
rect 2085 405 2143 439
rect 2085 371 2097 405
rect 2131 371 2143 405
rect 2085 355 2143 371
rect 2543 1629 2601 1645
rect 2543 1595 2555 1629
rect 2589 1595 2601 1629
rect 2543 1561 2601 1595
rect 2543 1527 2555 1561
rect 2589 1527 2601 1561
rect 2543 1493 2601 1527
rect 2543 1459 2555 1493
rect 2589 1459 2601 1493
rect 2543 1425 2601 1459
rect 2543 1391 2555 1425
rect 2589 1391 2601 1425
rect 2543 1357 2601 1391
rect 2543 1323 2555 1357
rect 2589 1323 2601 1357
rect 2543 1289 2601 1323
rect 2543 1255 2555 1289
rect 2589 1255 2601 1289
rect 2543 1221 2601 1255
rect 2543 1187 2555 1221
rect 2589 1187 2601 1221
rect 2543 1153 2601 1187
rect 2543 1119 2555 1153
rect 2589 1119 2601 1153
rect 2543 1085 2601 1119
rect 2543 1051 2555 1085
rect 2589 1051 2601 1085
rect 2543 1017 2601 1051
rect 2543 983 2555 1017
rect 2589 983 2601 1017
rect 2543 949 2601 983
rect 2543 915 2555 949
rect 2589 915 2601 949
rect 2543 881 2601 915
rect 2543 847 2555 881
rect 2589 847 2601 881
rect 2543 813 2601 847
rect 2543 779 2555 813
rect 2589 779 2601 813
rect 2543 745 2601 779
rect 2543 711 2555 745
rect 2589 711 2601 745
rect 2543 677 2601 711
rect 2543 643 2555 677
rect 2589 643 2601 677
rect 2543 609 2601 643
rect 2543 575 2555 609
rect 2589 575 2601 609
rect 2543 541 2601 575
rect 2543 507 2555 541
rect 2589 507 2601 541
rect 2543 473 2601 507
rect 2543 439 2555 473
rect 2589 439 2601 473
rect 2543 405 2601 439
rect 2543 371 2555 405
rect 2589 371 2601 405
rect 2543 355 2601 371
rect 3001 1629 3059 1645
rect 3001 1595 3013 1629
rect 3047 1595 3059 1629
rect 3001 1561 3059 1595
rect 3001 1527 3013 1561
rect 3047 1527 3059 1561
rect 3001 1493 3059 1527
rect 3001 1459 3013 1493
rect 3047 1459 3059 1493
rect 3001 1425 3059 1459
rect 3001 1391 3013 1425
rect 3047 1391 3059 1425
rect 3001 1357 3059 1391
rect 3001 1323 3013 1357
rect 3047 1323 3059 1357
rect 3001 1289 3059 1323
rect 3001 1255 3013 1289
rect 3047 1255 3059 1289
rect 3001 1221 3059 1255
rect 3001 1187 3013 1221
rect 3047 1187 3059 1221
rect 3001 1153 3059 1187
rect 3001 1119 3013 1153
rect 3047 1119 3059 1153
rect 3001 1085 3059 1119
rect 3001 1051 3013 1085
rect 3047 1051 3059 1085
rect 3001 1017 3059 1051
rect 3001 983 3013 1017
rect 3047 983 3059 1017
rect 3001 949 3059 983
rect 3001 915 3013 949
rect 3047 915 3059 949
rect 3001 881 3059 915
rect 3001 847 3013 881
rect 3047 847 3059 881
rect 3001 813 3059 847
rect 3001 779 3013 813
rect 3047 779 3059 813
rect 3001 745 3059 779
rect 3001 711 3013 745
rect 3047 711 3059 745
rect 3001 677 3059 711
rect 3001 643 3013 677
rect 3047 643 3059 677
rect 3001 609 3059 643
rect 3001 575 3013 609
rect 3047 575 3059 609
rect 3001 541 3059 575
rect 3001 507 3013 541
rect 3047 507 3059 541
rect 3001 473 3059 507
rect 3001 439 3013 473
rect 3047 439 3059 473
rect 3001 405 3059 439
rect 3001 371 3013 405
rect 3047 371 3059 405
rect 3001 355 3059 371
rect 3459 1629 3517 1645
rect 3459 1595 3471 1629
rect 3505 1595 3517 1629
rect 3459 1561 3517 1595
rect 3459 1527 3471 1561
rect 3505 1527 3517 1561
rect 3459 1493 3517 1527
rect 3459 1459 3471 1493
rect 3505 1459 3517 1493
rect 3459 1425 3517 1459
rect 3459 1391 3471 1425
rect 3505 1391 3517 1425
rect 3459 1357 3517 1391
rect 3459 1323 3471 1357
rect 3505 1323 3517 1357
rect 3459 1289 3517 1323
rect 3459 1255 3471 1289
rect 3505 1255 3517 1289
rect 3459 1221 3517 1255
rect 3459 1187 3471 1221
rect 3505 1187 3517 1221
rect 3459 1153 3517 1187
rect 3459 1119 3471 1153
rect 3505 1119 3517 1153
rect 3459 1085 3517 1119
rect 3459 1051 3471 1085
rect 3505 1051 3517 1085
rect 3459 1017 3517 1051
rect 3459 983 3471 1017
rect 3505 983 3517 1017
rect 3459 949 3517 983
rect 3459 915 3471 949
rect 3505 915 3517 949
rect 3459 881 3517 915
rect 3459 847 3471 881
rect 3505 847 3517 881
rect 3459 813 3517 847
rect 3459 779 3471 813
rect 3505 779 3517 813
rect 3459 745 3517 779
rect 3459 711 3471 745
rect 3505 711 3517 745
rect 3459 677 3517 711
rect 3459 643 3471 677
rect 3505 643 3517 677
rect 3459 609 3517 643
rect 3459 575 3471 609
rect 3505 575 3517 609
rect 3459 541 3517 575
rect 3459 507 3471 541
rect 3505 507 3517 541
rect 3459 473 3517 507
rect 3459 439 3471 473
rect 3505 439 3517 473
rect 3459 405 3517 439
rect 3459 371 3471 405
rect 3505 371 3517 405
rect 3459 355 3517 371
rect 3917 1629 3975 1645
rect 3917 1595 3929 1629
rect 3963 1595 3975 1629
rect 3917 1561 3975 1595
rect 3917 1527 3929 1561
rect 3963 1527 3975 1561
rect 3917 1493 3975 1527
rect 3917 1459 3929 1493
rect 3963 1459 3975 1493
rect 3917 1425 3975 1459
rect 3917 1391 3929 1425
rect 3963 1391 3975 1425
rect 3917 1357 3975 1391
rect 3917 1323 3929 1357
rect 3963 1323 3975 1357
rect 3917 1289 3975 1323
rect 3917 1255 3929 1289
rect 3963 1255 3975 1289
rect 3917 1221 3975 1255
rect 3917 1187 3929 1221
rect 3963 1187 3975 1221
rect 3917 1153 3975 1187
rect 3917 1119 3929 1153
rect 3963 1119 3975 1153
rect 3917 1085 3975 1119
rect 3917 1051 3929 1085
rect 3963 1051 3975 1085
rect 3917 1017 3975 1051
rect 3917 983 3929 1017
rect 3963 983 3975 1017
rect 3917 949 3975 983
rect 3917 915 3929 949
rect 3963 915 3975 949
rect 3917 881 3975 915
rect 3917 847 3929 881
rect 3963 847 3975 881
rect 3917 813 3975 847
rect 3917 779 3929 813
rect 3963 779 3975 813
rect 3917 745 3975 779
rect 3917 711 3929 745
rect 3963 711 3975 745
rect 3917 677 3975 711
rect 3917 643 3929 677
rect 3963 643 3975 677
rect 3917 609 3975 643
rect 3917 575 3929 609
rect 3963 575 3975 609
rect 3917 541 3975 575
rect 3917 507 3929 541
rect 3963 507 3975 541
rect 3917 473 3975 507
rect 3917 439 3929 473
rect 3963 439 3975 473
rect 3917 405 3975 439
rect 3917 371 3929 405
rect 3963 371 3975 405
rect 3917 355 3975 371
rect 4375 1629 4433 1645
rect 4375 1595 4387 1629
rect 4421 1595 4433 1629
rect 4375 1561 4433 1595
rect 4375 1527 4387 1561
rect 4421 1527 4433 1561
rect 4375 1493 4433 1527
rect 4375 1459 4387 1493
rect 4421 1459 4433 1493
rect 4375 1425 4433 1459
rect 4375 1391 4387 1425
rect 4421 1391 4433 1425
rect 4375 1357 4433 1391
rect 4375 1323 4387 1357
rect 4421 1323 4433 1357
rect 4375 1289 4433 1323
rect 4375 1255 4387 1289
rect 4421 1255 4433 1289
rect 4375 1221 4433 1255
rect 4375 1187 4387 1221
rect 4421 1187 4433 1221
rect 4375 1153 4433 1187
rect 4375 1119 4387 1153
rect 4421 1119 4433 1153
rect 4375 1085 4433 1119
rect 4375 1051 4387 1085
rect 4421 1051 4433 1085
rect 4375 1017 4433 1051
rect 4375 983 4387 1017
rect 4421 983 4433 1017
rect 4375 949 4433 983
rect 4375 915 4387 949
rect 4421 915 4433 949
rect 4375 881 4433 915
rect 4375 847 4387 881
rect 4421 847 4433 881
rect 4375 813 4433 847
rect 4375 779 4387 813
rect 4421 779 4433 813
rect 4375 745 4433 779
rect 4375 711 4387 745
rect 4421 711 4433 745
rect 4375 677 4433 711
rect 4375 643 4387 677
rect 4421 643 4433 677
rect 4375 609 4433 643
rect 4375 575 4387 609
rect 4421 575 4433 609
rect 4375 541 4433 575
rect 4375 507 4387 541
rect 4421 507 4433 541
rect 4375 473 4433 507
rect 4375 439 4387 473
rect 4421 439 4433 473
rect 4375 405 4433 439
rect 4375 371 4387 405
rect 4421 371 4433 405
rect 4375 355 4433 371
rect 4833 1629 4891 1645
rect 4833 1595 4845 1629
rect 4879 1595 4891 1629
rect 4833 1561 4891 1595
rect 4833 1527 4845 1561
rect 4879 1527 4891 1561
rect 4833 1493 4891 1527
rect 4833 1459 4845 1493
rect 4879 1459 4891 1493
rect 4833 1425 4891 1459
rect 4833 1391 4845 1425
rect 4879 1391 4891 1425
rect 4833 1357 4891 1391
rect 4833 1323 4845 1357
rect 4879 1323 4891 1357
rect 4833 1289 4891 1323
rect 4833 1255 4845 1289
rect 4879 1255 4891 1289
rect 4833 1221 4891 1255
rect 4833 1187 4845 1221
rect 4879 1187 4891 1221
rect 4833 1153 4891 1187
rect 4833 1119 4845 1153
rect 4879 1119 4891 1153
rect 4833 1085 4891 1119
rect 4833 1051 4845 1085
rect 4879 1051 4891 1085
rect 4833 1017 4891 1051
rect 4833 983 4845 1017
rect 4879 983 4891 1017
rect 4833 949 4891 983
rect 4833 915 4845 949
rect 4879 915 4891 949
rect 4833 881 4891 915
rect 4833 847 4845 881
rect 4879 847 4891 881
rect 4833 813 4891 847
rect 4833 779 4845 813
rect 4879 779 4891 813
rect 4833 745 4891 779
rect 4833 711 4845 745
rect 4879 711 4891 745
rect 4833 677 4891 711
rect 4833 643 4845 677
rect 4879 643 4891 677
rect 4833 609 4891 643
rect 4833 575 4845 609
rect 4879 575 4891 609
rect 4833 541 4891 575
rect 4833 507 4845 541
rect 4879 507 4891 541
rect 4833 473 4891 507
rect 4833 439 4845 473
rect 4879 439 4891 473
rect 4833 405 4891 439
rect 4833 371 4845 405
rect 4879 371 4891 405
rect 4833 355 4891 371
rect 5291 1629 5349 1645
rect 5291 1595 5303 1629
rect 5337 1595 5349 1629
rect 5291 1561 5349 1595
rect 5291 1527 5303 1561
rect 5337 1527 5349 1561
rect 5291 1493 5349 1527
rect 5291 1459 5303 1493
rect 5337 1459 5349 1493
rect 5291 1425 5349 1459
rect 5291 1391 5303 1425
rect 5337 1391 5349 1425
rect 5291 1357 5349 1391
rect 5291 1323 5303 1357
rect 5337 1323 5349 1357
rect 5291 1289 5349 1323
rect 5291 1255 5303 1289
rect 5337 1255 5349 1289
rect 5291 1221 5349 1255
rect 5291 1187 5303 1221
rect 5337 1187 5349 1221
rect 5291 1153 5349 1187
rect 5291 1119 5303 1153
rect 5337 1119 5349 1153
rect 5291 1085 5349 1119
rect 5291 1051 5303 1085
rect 5337 1051 5349 1085
rect 5291 1017 5349 1051
rect 5291 983 5303 1017
rect 5337 983 5349 1017
rect 5291 949 5349 983
rect 5291 915 5303 949
rect 5337 915 5349 949
rect 5291 881 5349 915
rect 5291 847 5303 881
rect 5337 847 5349 881
rect 5291 813 5349 847
rect 5291 779 5303 813
rect 5337 779 5349 813
rect 5291 745 5349 779
rect 5291 711 5303 745
rect 5337 711 5349 745
rect 5291 677 5349 711
rect 5291 643 5303 677
rect 5337 643 5349 677
rect 5291 609 5349 643
rect 5291 575 5303 609
rect 5337 575 5349 609
rect 5291 541 5349 575
rect 5291 507 5303 541
rect 5337 507 5349 541
rect 5291 473 5349 507
rect 5291 439 5303 473
rect 5337 439 5349 473
rect 5291 405 5349 439
rect 5291 371 5303 405
rect 5337 371 5349 405
rect 5291 355 5349 371
rect 5749 1629 5807 1645
rect 5749 1595 5761 1629
rect 5795 1595 5807 1629
rect 5749 1561 5807 1595
rect 5749 1527 5761 1561
rect 5795 1527 5807 1561
rect 5749 1493 5807 1527
rect 5749 1459 5761 1493
rect 5795 1459 5807 1493
rect 5749 1425 5807 1459
rect 5749 1391 5761 1425
rect 5795 1391 5807 1425
rect 5749 1357 5807 1391
rect 5749 1323 5761 1357
rect 5795 1323 5807 1357
rect 5749 1289 5807 1323
rect 5749 1255 5761 1289
rect 5795 1255 5807 1289
rect 5749 1221 5807 1255
rect 5749 1187 5761 1221
rect 5795 1187 5807 1221
rect 5749 1153 5807 1187
rect 5749 1119 5761 1153
rect 5795 1119 5807 1153
rect 5749 1085 5807 1119
rect 5749 1051 5761 1085
rect 5795 1051 5807 1085
rect 5749 1017 5807 1051
rect 5749 983 5761 1017
rect 5795 983 5807 1017
rect 5749 949 5807 983
rect 5749 915 5761 949
rect 5795 915 5807 949
rect 5749 881 5807 915
rect 5749 847 5761 881
rect 5795 847 5807 881
rect 5749 813 5807 847
rect 5749 779 5761 813
rect 5795 779 5807 813
rect 5749 745 5807 779
rect 5749 711 5761 745
rect 5795 711 5807 745
rect 5749 677 5807 711
rect 5749 643 5761 677
rect 5795 643 5807 677
rect 5749 609 5807 643
rect 5749 575 5761 609
rect 5795 575 5807 609
rect 5749 541 5807 575
rect 5749 507 5761 541
rect 5795 507 5807 541
rect 5749 473 5807 507
rect 5749 439 5761 473
rect 5795 439 5807 473
rect 5749 405 5807 439
rect 5749 371 5761 405
rect 5795 371 5807 405
rect 5749 355 5807 371
<< pdiffc >>
rect 265 1595 299 1629
rect 265 1527 299 1561
rect 265 1459 299 1493
rect 265 1391 299 1425
rect 265 1323 299 1357
rect 265 1255 299 1289
rect 265 1187 299 1221
rect 265 1119 299 1153
rect 265 1051 299 1085
rect 265 983 299 1017
rect 265 915 299 949
rect 265 847 299 881
rect 265 779 299 813
rect 265 711 299 745
rect 265 643 299 677
rect 265 575 299 609
rect 265 507 299 541
rect 265 439 299 473
rect 265 371 299 405
rect 723 1595 757 1629
rect 723 1527 757 1561
rect 723 1459 757 1493
rect 723 1391 757 1425
rect 723 1323 757 1357
rect 723 1255 757 1289
rect 723 1187 757 1221
rect 723 1119 757 1153
rect 723 1051 757 1085
rect 723 983 757 1017
rect 723 915 757 949
rect 723 847 757 881
rect 723 779 757 813
rect 723 711 757 745
rect 723 643 757 677
rect 723 575 757 609
rect 723 507 757 541
rect 723 439 757 473
rect 723 371 757 405
rect 1181 1595 1215 1629
rect 1181 1527 1215 1561
rect 1181 1459 1215 1493
rect 1181 1391 1215 1425
rect 1181 1323 1215 1357
rect 1181 1255 1215 1289
rect 1181 1187 1215 1221
rect 1181 1119 1215 1153
rect 1181 1051 1215 1085
rect 1181 983 1215 1017
rect 1181 915 1215 949
rect 1181 847 1215 881
rect 1181 779 1215 813
rect 1181 711 1215 745
rect 1181 643 1215 677
rect 1181 575 1215 609
rect 1181 507 1215 541
rect 1181 439 1215 473
rect 1181 371 1215 405
rect 1639 1595 1673 1629
rect 1639 1527 1673 1561
rect 1639 1459 1673 1493
rect 1639 1391 1673 1425
rect 1639 1323 1673 1357
rect 1639 1255 1673 1289
rect 1639 1187 1673 1221
rect 1639 1119 1673 1153
rect 1639 1051 1673 1085
rect 1639 983 1673 1017
rect 1639 915 1673 949
rect 1639 847 1673 881
rect 1639 779 1673 813
rect 1639 711 1673 745
rect 1639 643 1673 677
rect 1639 575 1673 609
rect 1639 507 1673 541
rect 1639 439 1673 473
rect 1639 371 1673 405
rect 2097 1595 2131 1629
rect 2097 1527 2131 1561
rect 2097 1459 2131 1493
rect 2097 1391 2131 1425
rect 2097 1323 2131 1357
rect 2097 1255 2131 1289
rect 2097 1187 2131 1221
rect 2097 1119 2131 1153
rect 2097 1051 2131 1085
rect 2097 983 2131 1017
rect 2097 915 2131 949
rect 2097 847 2131 881
rect 2097 779 2131 813
rect 2097 711 2131 745
rect 2097 643 2131 677
rect 2097 575 2131 609
rect 2097 507 2131 541
rect 2097 439 2131 473
rect 2097 371 2131 405
rect 2555 1595 2589 1629
rect 2555 1527 2589 1561
rect 2555 1459 2589 1493
rect 2555 1391 2589 1425
rect 2555 1323 2589 1357
rect 2555 1255 2589 1289
rect 2555 1187 2589 1221
rect 2555 1119 2589 1153
rect 2555 1051 2589 1085
rect 2555 983 2589 1017
rect 2555 915 2589 949
rect 2555 847 2589 881
rect 2555 779 2589 813
rect 2555 711 2589 745
rect 2555 643 2589 677
rect 2555 575 2589 609
rect 2555 507 2589 541
rect 2555 439 2589 473
rect 2555 371 2589 405
rect 3013 1595 3047 1629
rect 3013 1527 3047 1561
rect 3013 1459 3047 1493
rect 3013 1391 3047 1425
rect 3013 1323 3047 1357
rect 3013 1255 3047 1289
rect 3013 1187 3047 1221
rect 3013 1119 3047 1153
rect 3013 1051 3047 1085
rect 3013 983 3047 1017
rect 3013 915 3047 949
rect 3013 847 3047 881
rect 3013 779 3047 813
rect 3013 711 3047 745
rect 3013 643 3047 677
rect 3013 575 3047 609
rect 3013 507 3047 541
rect 3013 439 3047 473
rect 3013 371 3047 405
rect 3471 1595 3505 1629
rect 3471 1527 3505 1561
rect 3471 1459 3505 1493
rect 3471 1391 3505 1425
rect 3471 1323 3505 1357
rect 3471 1255 3505 1289
rect 3471 1187 3505 1221
rect 3471 1119 3505 1153
rect 3471 1051 3505 1085
rect 3471 983 3505 1017
rect 3471 915 3505 949
rect 3471 847 3505 881
rect 3471 779 3505 813
rect 3471 711 3505 745
rect 3471 643 3505 677
rect 3471 575 3505 609
rect 3471 507 3505 541
rect 3471 439 3505 473
rect 3471 371 3505 405
rect 3929 1595 3963 1629
rect 3929 1527 3963 1561
rect 3929 1459 3963 1493
rect 3929 1391 3963 1425
rect 3929 1323 3963 1357
rect 3929 1255 3963 1289
rect 3929 1187 3963 1221
rect 3929 1119 3963 1153
rect 3929 1051 3963 1085
rect 3929 983 3963 1017
rect 3929 915 3963 949
rect 3929 847 3963 881
rect 3929 779 3963 813
rect 3929 711 3963 745
rect 3929 643 3963 677
rect 3929 575 3963 609
rect 3929 507 3963 541
rect 3929 439 3963 473
rect 3929 371 3963 405
rect 4387 1595 4421 1629
rect 4387 1527 4421 1561
rect 4387 1459 4421 1493
rect 4387 1391 4421 1425
rect 4387 1323 4421 1357
rect 4387 1255 4421 1289
rect 4387 1187 4421 1221
rect 4387 1119 4421 1153
rect 4387 1051 4421 1085
rect 4387 983 4421 1017
rect 4387 915 4421 949
rect 4387 847 4421 881
rect 4387 779 4421 813
rect 4387 711 4421 745
rect 4387 643 4421 677
rect 4387 575 4421 609
rect 4387 507 4421 541
rect 4387 439 4421 473
rect 4387 371 4421 405
rect 4845 1595 4879 1629
rect 4845 1527 4879 1561
rect 4845 1459 4879 1493
rect 4845 1391 4879 1425
rect 4845 1323 4879 1357
rect 4845 1255 4879 1289
rect 4845 1187 4879 1221
rect 4845 1119 4879 1153
rect 4845 1051 4879 1085
rect 4845 983 4879 1017
rect 4845 915 4879 949
rect 4845 847 4879 881
rect 4845 779 4879 813
rect 4845 711 4879 745
rect 4845 643 4879 677
rect 4845 575 4879 609
rect 4845 507 4879 541
rect 4845 439 4879 473
rect 4845 371 4879 405
rect 5303 1595 5337 1629
rect 5303 1527 5337 1561
rect 5303 1459 5337 1493
rect 5303 1391 5337 1425
rect 5303 1323 5337 1357
rect 5303 1255 5337 1289
rect 5303 1187 5337 1221
rect 5303 1119 5337 1153
rect 5303 1051 5337 1085
rect 5303 983 5337 1017
rect 5303 915 5337 949
rect 5303 847 5337 881
rect 5303 779 5337 813
rect 5303 711 5337 745
rect 5303 643 5337 677
rect 5303 575 5337 609
rect 5303 507 5337 541
rect 5303 439 5337 473
rect 5303 371 5337 405
rect 5761 1595 5795 1629
rect 5761 1527 5795 1561
rect 5761 1459 5795 1493
rect 5761 1391 5795 1425
rect 5761 1323 5795 1357
rect 5761 1255 5795 1289
rect 5761 1187 5795 1221
rect 5761 1119 5795 1153
rect 5761 1051 5795 1085
rect 5761 983 5795 1017
rect 5761 915 5795 949
rect 5761 847 5795 881
rect 5761 779 5795 813
rect 5761 711 5795 745
rect 5761 643 5795 677
rect 5761 575 5795 609
rect 5761 507 5795 541
rect 5761 439 5795 473
rect 5761 371 5795 405
<< nsubdiff >>
rect 1216 1807 1336 1810
rect 158 1757 198 1800
rect 1216 1773 1261 1807
rect 1295 1773 1336 1807
rect 1216 1770 1336 1773
rect 2516 1807 2636 1810
rect 2516 1773 2561 1807
rect 2595 1773 2636 1807
rect 2516 1770 2636 1773
rect 3816 1807 3936 1810
rect 3816 1773 3861 1807
rect 3895 1773 3936 1807
rect 3816 1770 3936 1773
rect 158 1723 161 1757
rect 195 1723 198 1757
rect 158 1680 198 1723
<< nsubdiffcont >>
rect 1261 1773 1295 1807
rect 2561 1773 2595 1807
rect 3861 1773 3895 1807
rect 161 1723 195 1757
<< poly >>
rect 311 1645 711 1671
rect 769 1645 1169 1671
rect 1227 1645 1627 1671
rect 1685 1645 2085 1671
rect 2143 1645 2543 1671
rect 2601 1645 3001 1671
rect 3059 1645 3459 1671
rect 3517 1645 3917 1671
rect 3975 1645 4375 1671
rect 4433 1645 4833 1671
rect 4891 1645 5291 1671
rect 5349 1645 5749 1671
rect 311 329 711 355
rect 769 329 1169 355
rect 1227 329 1627 355
rect 1685 329 2085 355
rect 2143 329 2543 355
rect 2601 329 3001 355
rect 3059 329 3459 355
rect 3517 329 3917 355
rect 3975 329 4375 355
rect 4433 329 4833 355
rect 4891 329 5291 355
rect 5349 329 5749 355
rect 458 184 578 329
rect 914 184 1034 329
rect 1370 184 1490 329
rect 1826 184 1946 329
rect 2282 184 2402 329
rect 2738 184 2858 329
rect 3194 184 3314 329
rect 3650 184 3770 329
rect 4106 184 4226 329
rect 4562 184 4682 329
rect 5018 184 5138 329
rect 5474 184 5594 329
rect 218 151 5842 184
rect 218 117 401 151
rect 435 117 801 151
rect 835 117 1201 151
rect 1235 117 1601 151
rect 1635 117 2001 151
rect 2035 117 2401 151
rect 2435 117 2801 151
rect 2835 117 3201 151
rect 3235 117 3601 151
rect 3635 117 4001 151
rect 4035 117 4401 151
rect 4435 117 4801 151
rect 4835 117 5201 151
rect 5235 117 5601 151
rect 5635 117 5842 151
rect 218 84 5842 117
<< polycont >>
rect 401 117 435 151
rect 801 117 835 151
rect 1201 117 1235 151
rect 1601 117 1635 151
rect 2001 117 2035 151
rect 2401 117 2435 151
rect 2801 117 2835 151
rect 3201 117 3235 151
rect 3601 117 3635 151
rect 4001 117 4035 151
rect 4401 117 4435 151
rect 4801 117 4835 151
rect 5201 117 5235 151
rect 5601 117 5635 151
<< locali >>
rect 120 1897 5842 1910
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3201 1897
rect 3235 1863 3601 1897
rect 3635 1863 4001 1897
rect 4035 1863 4401 1897
rect 4435 1863 4801 1897
rect 4835 1863 5201 1897
rect 5235 1863 5601 1897
rect 5635 1863 5842 1897
rect 120 1850 5842 1863
rect 148 1757 208 1850
rect 1196 1807 1356 1850
rect 1196 1773 1261 1807
rect 1295 1773 1356 1807
rect 1196 1770 1356 1773
rect 2496 1807 2656 1850
rect 2496 1773 2561 1807
rect 2595 1773 2656 1807
rect 2496 1770 2656 1773
rect 3796 1807 3956 1850
rect 3796 1773 3861 1807
rect 3895 1773 3956 1807
rect 3796 1770 3956 1773
rect 148 1723 161 1757
rect 195 1723 208 1757
rect 148 1640 208 1723
rect 278 1690 5842 1730
rect 265 1629 299 1649
rect 265 1561 299 1595
rect 265 1493 299 1523
rect 265 1425 299 1451
rect 265 1357 299 1379
rect 265 1289 299 1307
rect 265 1221 299 1235
rect 265 1153 299 1163
rect 265 1085 299 1091
rect 265 1017 299 1019
rect 265 981 299 983
rect 265 909 299 915
rect 265 837 299 847
rect 265 765 299 779
rect 265 693 299 711
rect 265 621 299 643
rect 265 549 299 575
rect 265 477 299 507
rect 265 405 299 439
rect 265 270 299 371
rect 723 1629 757 1690
rect 723 1561 757 1595
rect 723 1493 757 1523
rect 723 1425 757 1451
rect 723 1357 757 1379
rect 723 1289 757 1307
rect 723 1221 757 1235
rect 723 1153 757 1163
rect 723 1085 757 1091
rect 723 1017 757 1019
rect 723 981 757 983
rect 723 909 757 915
rect 723 837 757 847
rect 723 765 757 779
rect 723 693 757 711
rect 723 621 757 643
rect 723 549 757 575
rect 723 477 757 507
rect 723 405 757 439
rect 723 351 757 371
rect 1181 1629 1215 1649
rect 1181 1561 1215 1595
rect 1181 1493 1215 1523
rect 1181 1425 1215 1451
rect 1181 1357 1215 1379
rect 1181 1289 1215 1307
rect 1181 1221 1215 1235
rect 1181 1153 1215 1163
rect 1181 1085 1215 1091
rect 1181 1017 1215 1019
rect 1181 981 1215 983
rect 1181 909 1215 915
rect 1181 837 1215 847
rect 1181 765 1215 779
rect 1181 693 1215 711
rect 1181 621 1215 643
rect 1181 549 1215 575
rect 1181 477 1215 507
rect 1181 405 1215 439
rect 1181 270 1215 371
rect 1639 1629 1673 1690
rect 1639 1561 1673 1595
rect 1639 1493 1673 1523
rect 1639 1425 1673 1451
rect 1639 1357 1673 1379
rect 1639 1289 1673 1307
rect 1639 1221 1673 1235
rect 1639 1153 1673 1163
rect 1639 1085 1673 1091
rect 1639 1017 1673 1019
rect 1639 981 1673 983
rect 1639 909 1673 915
rect 1639 837 1673 847
rect 1639 765 1673 779
rect 1639 693 1673 711
rect 1639 621 1673 643
rect 1639 549 1673 575
rect 1639 477 1673 507
rect 1639 405 1673 439
rect 1639 351 1673 371
rect 2097 1629 2131 1649
rect 2097 1561 2131 1595
rect 2097 1493 2131 1523
rect 2097 1425 2131 1451
rect 2097 1357 2131 1379
rect 2097 1289 2131 1307
rect 2097 1221 2131 1235
rect 2097 1153 2131 1163
rect 2097 1085 2131 1091
rect 2097 1017 2131 1019
rect 2097 981 2131 983
rect 2097 909 2131 915
rect 2097 837 2131 847
rect 2097 765 2131 779
rect 2097 693 2131 711
rect 2097 621 2131 643
rect 2097 549 2131 575
rect 2097 477 2131 507
rect 2097 405 2131 439
rect 2097 270 2131 371
rect 2555 1629 2589 1690
rect 2555 1561 2589 1595
rect 2555 1493 2589 1523
rect 2555 1425 2589 1451
rect 2555 1357 2589 1379
rect 2555 1289 2589 1307
rect 2555 1221 2589 1235
rect 2555 1153 2589 1163
rect 2555 1085 2589 1091
rect 2555 1017 2589 1019
rect 2555 981 2589 983
rect 2555 909 2589 915
rect 2555 837 2589 847
rect 2555 765 2589 779
rect 2555 693 2589 711
rect 2555 621 2589 643
rect 2555 549 2589 575
rect 2555 477 2589 507
rect 2555 405 2589 439
rect 2555 351 2589 371
rect 3013 1629 3047 1649
rect 3013 1561 3047 1595
rect 3013 1493 3047 1523
rect 3013 1425 3047 1451
rect 3013 1357 3047 1379
rect 3013 1289 3047 1307
rect 3013 1221 3047 1235
rect 3013 1153 3047 1163
rect 3013 1085 3047 1091
rect 3013 1017 3047 1019
rect 3013 981 3047 983
rect 3013 909 3047 915
rect 3013 837 3047 847
rect 3013 765 3047 779
rect 3013 693 3047 711
rect 3013 621 3047 643
rect 3013 549 3047 575
rect 3013 477 3047 507
rect 3013 405 3047 439
rect 3013 270 3047 371
rect 3471 1629 3505 1690
rect 3471 1561 3505 1595
rect 3471 1493 3505 1523
rect 3471 1425 3505 1451
rect 3471 1357 3505 1379
rect 3471 1289 3505 1307
rect 3471 1221 3505 1235
rect 3471 1153 3505 1163
rect 3471 1085 3505 1091
rect 3471 1017 3505 1019
rect 3471 981 3505 983
rect 3471 909 3505 915
rect 3471 837 3505 847
rect 3471 765 3505 779
rect 3471 693 3505 711
rect 3471 621 3505 643
rect 3471 549 3505 575
rect 3471 477 3505 507
rect 3471 405 3505 439
rect 3471 351 3505 371
rect 3929 1629 3963 1649
rect 3929 1561 3963 1595
rect 3929 1493 3963 1523
rect 3929 1425 3963 1451
rect 3929 1357 3963 1379
rect 3929 1289 3963 1307
rect 3929 1221 3963 1235
rect 3929 1153 3963 1163
rect 3929 1085 3963 1091
rect 3929 1017 3963 1019
rect 3929 981 3963 983
rect 3929 909 3963 915
rect 3929 837 3963 847
rect 3929 765 3963 779
rect 3929 693 3963 711
rect 3929 621 3963 643
rect 3929 549 3963 575
rect 3929 477 3963 507
rect 3929 405 3963 439
rect 3929 270 3963 371
rect 4387 1629 4421 1690
rect 4387 1561 4421 1595
rect 4387 1493 4421 1523
rect 4387 1425 4421 1451
rect 4387 1357 4421 1379
rect 4387 1289 4421 1307
rect 4387 1221 4421 1235
rect 4387 1153 4421 1163
rect 4387 1085 4421 1091
rect 4387 1017 4421 1019
rect 4387 981 4421 983
rect 4387 909 4421 915
rect 4387 837 4421 847
rect 4387 765 4421 779
rect 4387 693 4421 711
rect 4387 621 4421 643
rect 4387 549 4421 575
rect 4387 477 4421 507
rect 4387 405 4421 439
rect 4387 351 4421 371
rect 4845 1629 4879 1649
rect 4845 1561 4879 1595
rect 4845 1493 4879 1523
rect 4845 1425 4879 1451
rect 4845 1357 4879 1379
rect 4845 1289 4879 1307
rect 4845 1221 4879 1235
rect 4845 1153 4879 1163
rect 4845 1085 4879 1091
rect 4845 1017 4879 1019
rect 4845 981 4879 983
rect 4845 909 4879 915
rect 4845 837 4879 847
rect 4845 765 4879 779
rect 4845 693 4879 711
rect 4845 621 4879 643
rect 4845 549 4879 575
rect 4845 477 4879 507
rect 4845 405 4879 439
rect 4845 270 4879 371
rect 5303 1629 5337 1690
rect 5303 1561 5337 1595
rect 5303 1493 5337 1523
rect 5303 1425 5337 1451
rect 5303 1357 5337 1379
rect 5303 1289 5337 1307
rect 5303 1221 5337 1235
rect 5303 1153 5337 1163
rect 5303 1085 5337 1091
rect 5303 1017 5337 1019
rect 5303 981 5337 983
rect 5303 909 5337 915
rect 5303 837 5337 847
rect 5303 765 5337 779
rect 5303 693 5337 711
rect 5303 621 5337 643
rect 5303 549 5337 575
rect 5303 477 5337 507
rect 5303 405 5337 439
rect 5303 351 5337 371
rect 5761 1629 5795 1649
rect 5761 1561 5795 1595
rect 5761 1493 5795 1523
rect 5761 1425 5795 1451
rect 5761 1357 5795 1379
rect 5761 1289 5795 1307
rect 5761 1221 5795 1235
rect 5761 1153 5795 1163
rect 5761 1085 5795 1091
rect 5761 1017 5795 1019
rect 5761 981 5795 983
rect 5761 909 5795 915
rect 5761 837 5795 847
rect 5761 765 5795 779
rect 5761 693 5795 711
rect 5761 621 5795 643
rect 5761 549 5795 575
rect 5761 477 5795 507
rect 5761 405 5795 439
rect 5761 270 5795 371
rect 218 210 5842 270
rect 218 151 5842 164
rect 218 117 401 151
rect 435 117 801 151
rect 835 117 1201 151
rect 1235 117 1601 151
rect 1635 117 2001 151
rect 2035 117 2401 151
rect 2435 117 2801 151
rect 2835 117 3201 151
rect 3235 117 3601 151
rect 3635 117 4001 151
rect 4035 117 4401 151
rect 4435 117 4801 151
rect 4835 117 5201 151
rect 5235 117 5601 151
rect 5635 117 5842 151
rect 218 104 5842 117
rect 120 17 5842 30
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3201 17
rect 3235 -17 3601 17
rect 3635 -17 4001 17
rect 4035 -17 4401 17
rect 4435 -17 4801 17
rect 4835 -17 5201 17
rect 5235 -17 5601 17
rect 5635 -17 5842 17
rect 120 -30 5842 -17
<< viali >>
rect 401 1863 435 1897
rect 801 1863 835 1897
rect 1201 1863 1235 1897
rect 1601 1863 1635 1897
rect 2001 1863 2035 1897
rect 2401 1863 2435 1897
rect 2801 1863 2835 1897
rect 3201 1863 3235 1897
rect 3601 1863 3635 1897
rect 4001 1863 4035 1897
rect 4401 1863 4435 1897
rect 4801 1863 4835 1897
rect 5201 1863 5235 1897
rect 5601 1863 5635 1897
rect 265 1595 299 1629
rect 265 1527 299 1557
rect 265 1523 299 1527
rect 265 1459 299 1485
rect 265 1451 299 1459
rect 265 1391 299 1413
rect 265 1379 299 1391
rect 265 1323 299 1341
rect 265 1307 299 1323
rect 265 1255 299 1269
rect 265 1235 299 1255
rect 265 1187 299 1197
rect 265 1163 299 1187
rect 265 1119 299 1125
rect 265 1091 299 1119
rect 265 1051 299 1053
rect 265 1019 299 1051
rect 265 949 299 981
rect 265 947 299 949
rect 265 881 299 909
rect 265 875 299 881
rect 265 813 299 837
rect 265 803 299 813
rect 265 745 299 765
rect 265 731 299 745
rect 265 677 299 693
rect 265 659 299 677
rect 265 609 299 621
rect 265 587 299 609
rect 265 541 299 549
rect 265 515 299 541
rect 265 473 299 477
rect 265 443 299 473
rect 265 371 299 405
rect 723 1595 757 1629
rect 723 1527 757 1557
rect 723 1523 757 1527
rect 723 1459 757 1485
rect 723 1451 757 1459
rect 723 1391 757 1413
rect 723 1379 757 1391
rect 723 1323 757 1341
rect 723 1307 757 1323
rect 723 1255 757 1269
rect 723 1235 757 1255
rect 723 1187 757 1197
rect 723 1163 757 1187
rect 723 1119 757 1125
rect 723 1091 757 1119
rect 723 1051 757 1053
rect 723 1019 757 1051
rect 723 949 757 981
rect 723 947 757 949
rect 723 881 757 909
rect 723 875 757 881
rect 723 813 757 837
rect 723 803 757 813
rect 723 745 757 765
rect 723 731 757 745
rect 723 677 757 693
rect 723 659 757 677
rect 723 609 757 621
rect 723 587 757 609
rect 723 541 757 549
rect 723 515 757 541
rect 723 473 757 477
rect 723 443 757 473
rect 723 371 757 405
rect 1181 1595 1215 1629
rect 1181 1527 1215 1557
rect 1181 1523 1215 1527
rect 1181 1459 1215 1485
rect 1181 1451 1215 1459
rect 1181 1391 1215 1413
rect 1181 1379 1215 1391
rect 1181 1323 1215 1341
rect 1181 1307 1215 1323
rect 1181 1255 1215 1269
rect 1181 1235 1215 1255
rect 1181 1187 1215 1197
rect 1181 1163 1215 1187
rect 1181 1119 1215 1125
rect 1181 1091 1215 1119
rect 1181 1051 1215 1053
rect 1181 1019 1215 1051
rect 1181 949 1215 981
rect 1181 947 1215 949
rect 1181 881 1215 909
rect 1181 875 1215 881
rect 1181 813 1215 837
rect 1181 803 1215 813
rect 1181 745 1215 765
rect 1181 731 1215 745
rect 1181 677 1215 693
rect 1181 659 1215 677
rect 1181 609 1215 621
rect 1181 587 1215 609
rect 1181 541 1215 549
rect 1181 515 1215 541
rect 1181 473 1215 477
rect 1181 443 1215 473
rect 1181 371 1215 405
rect 1639 1595 1673 1629
rect 1639 1527 1673 1557
rect 1639 1523 1673 1527
rect 1639 1459 1673 1485
rect 1639 1451 1673 1459
rect 1639 1391 1673 1413
rect 1639 1379 1673 1391
rect 1639 1323 1673 1341
rect 1639 1307 1673 1323
rect 1639 1255 1673 1269
rect 1639 1235 1673 1255
rect 1639 1187 1673 1197
rect 1639 1163 1673 1187
rect 1639 1119 1673 1125
rect 1639 1091 1673 1119
rect 1639 1051 1673 1053
rect 1639 1019 1673 1051
rect 1639 949 1673 981
rect 1639 947 1673 949
rect 1639 881 1673 909
rect 1639 875 1673 881
rect 1639 813 1673 837
rect 1639 803 1673 813
rect 1639 745 1673 765
rect 1639 731 1673 745
rect 1639 677 1673 693
rect 1639 659 1673 677
rect 1639 609 1673 621
rect 1639 587 1673 609
rect 1639 541 1673 549
rect 1639 515 1673 541
rect 1639 473 1673 477
rect 1639 443 1673 473
rect 1639 371 1673 405
rect 2097 1595 2131 1629
rect 2097 1527 2131 1557
rect 2097 1523 2131 1527
rect 2097 1459 2131 1485
rect 2097 1451 2131 1459
rect 2097 1391 2131 1413
rect 2097 1379 2131 1391
rect 2097 1323 2131 1341
rect 2097 1307 2131 1323
rect 2097 1255 2131 1269
rect 2097 1235 2131 1255
rect 2097 1187 2131 1197
rect 2097 1163 2131 1187
rect 2097 1119 2131 1125
rect 2097 1091 2131 1119
rect 2097 1051 2131 1053
rect 2097 1019 2131 1051
rect 2097 949 2131 981
rect 2097 947 2131 949
rect 2097 881 2131 909
rect 2097 875 2131 881
rect 2097 813 2131 837
rect 2097 803 2131 813
rect 2097 745 2131 765
rect 2097 731 2131 745
rect 2097 677 2131 693
rect 2097 659 2131 677
rect 2097 609 2131 621
rect 2097 587 2131 609
rect 2097 541 2131 549
rect 2097 515 2131 541
rect 2097 473 2131 477
rect 2097 443 2131 473
rect 2097 371 2131 405
rect 2555 1595 2589 1629
rect 2555 1527 2589 1557
rect 2555 1523 2589 1527
rect 2555 1459 2589 1485
rect 2555 1451 2589 1459
rect 2555 1391 2589 1413
rect 2555 1379 2589 1391
rect 2555 1323 2589 1341
rect 2555 1307 2589 1323
rect 2555 1255 2589 1269
rect 2555 1235 2589 1255
rect 2555 1187 2589 1197
rect 2555 1163 2589 1187
rect 2555 1119 2589 1125
rect 2555 1091 2589 1119
rect 2555 1051 2589 1053
rect 2555 1019 2589 1051
rect 2555 949 2589 981
rect 2555 947 2589 949
rect 2555 881 2589 909
rect 2555 875 2589 881
rect 2555 813 2589 837
rect 2555 803 2589 813
rect 2555 745 2589 765
rect 2555 731 2589 745
rect 2555 677 2589 693
rect 2555 659 2589 677
rect 2555 609 2589 621
rect 2555 587 2589 609
rect 2555 541 2589 549
rect 2555 515 2589 541
rect 2555 473 2589 477
rect 2555 443 2589 473
rect 2555 371 2589 405
rect 3013 1595 3047 1629
rect 3013 1527 3047 1557
rect 3013 1523 3047 1527
rect 3013 1459 3047 1485
rect 3013 1451 3047 1459
rect 3013 1391 3047 1413
rect 3013 1379 3047 1391
rect 3013 1323 3047 1341
rect 3013 1307 3047 1323
rect 3013 1255 3047 1269
rect 3013 1235 3047 1255
rect 3013 1187 3047 1197
rect 3013 1163 3047 1187
rect 3013 1119 3047 1125
rect 3013 1091 3047 1119
rect 3013 1051 3047 1053
rect 3013 1019 3047 1051
rect 3013 949 3047 981
rect 3013 947 3047 949
rect 3013 881 3047 909
rect 3013 875 3047 881
rect 3013 813 3047 837
rect 3013 803 3047 813
rect 3013 745 3047 765
rect 3013 731 3047 745
rect 3013 677 3047 693
rect 3013 659 3047 677
rect 3013 609 3047 621
rect 3013 587 3047 609
rect 3013 541 3047 549
rect 3013 515 3047 541
rect 3013 473 3047 477
rect 3013 443 3047 473
rect 3013 371 3047 405
rect 3471 1595 3505 1629
rect 3471 1527 3505 1557
rect 3471 1523 3505 1527
rect 3471 1459 3505 1485
rect 3471 1451 3505 1459
rect 3471 1391 3505 1413
rect 3471 1379 3505 1391
rect 3471 1323 3505 1341
rect 3471 1307 3505 1323
rect 3471 1255 3505 1269
rect 3471 1235 3505 1255
rect 3471 1187 3505 1197
rect 3471 1163 3505 1187
rect 3471 1119 3505 1125
rect 3471 1091 3505 1119
rect 3471 1051 3505 1053
rect 3471 1019 3505 1051
rect 3471 949 3505 981
rect 3471 947 3505 949
rect 3471 881 3505 909
rect 3471 875 3505 881
rect 3471 813 3505 837
rect 3471 803 3505 813
rect 3471 745 3505 765
rect 3471 731 3505 745
rect 3471 677 3505 693
rect 3471 659 3505 677
rect 3471 609 3505 621
rect 3471 587 3505 609
rect 3471 541 3505 549
rect 3471 515 3505 541
rect 3471 473 3505 477
rect 3471 443 3505 473
rect 3471 371 3505 405
rect 3929 1595 3963 1629
rect 3929 1527 3963 1557
rect 3929 1523 3963 1527
rect 3929 1459 3963 1485
rect 3929 1451 3963 1459
rect 3929 1391 3963 1413
rect 3929 1379 3963 1391
rect 3929 1323 3963 1341
rect 3929 1307 3963 1323
rect 3929 1255 3963 1269
rect 3929 1235 3963 1255
rect 3929 1187 3963 1197
rect 3929 1163 3963 1187
rect 3929 1119 3963 1125
rect 3929 1091 3963 1119
rect 3929 1051 3963 1053
rect 3929 1019 3963 1051
rect 3929 949 3963 981
rect 3929 947 3963 949
rect 3929 881 3963 909
rect 3929 875 3963 881
rect 3929 813 3963 837
rect 3929 803 3963 813
rect 3929 745 3963 765
rect 3929 731 3963 745
rect 3929 677 3963 693
rect 3929 659 3963 677
rect 3929 609 3963 621
rect 3929 587 3963 609
rect 3929 541 3963 549
rect 3929 515 3963 541
rect 3929 473 3963 477
rect 3929 443 3963 473
rect 3929 371 3963 405
rect 4387 1595 4421 1629
rect 4387 1527 4421 1557
rect 4387 1523 4421 1527
rect 4387 1459 4421 1485
rect 4387 1451 4421 1459
rect 4387 1391 4421 1413
rect 4387 1379 4421 1391
rect 4387 1323 4421 1341
rect 4387 1307 4421 1323
rect 4387 1255 4421 1269
rect 4387 1235 4421 1255
rect 4387 1187 4421 1197
rect 4387 1163 4421 1187
rect 4387 1119 4421 1125
rect 4387 1091 4421 1119
rect 4387 1051 4421 1053
rect 4387 1019 4421 1051
rect 4387 949 4421 981
rect 4387 947 4421 949
rect 4387 881 4421 909
rect 4387 875 4421 881
rect 4387 813 4421 837
rect 4387 803 4421 813
rect 4387 745 4421 765
rect 4387 731 4421 745
rect 4387 677 4421 693
rect 4387 659 4421 677
rect 4387 609 4421 621
rect 4387 587 4421 609
rect 4387 541 4421 549
rect 4387 515 4421 541
rect 4387 473 4421 477
rect 4387 443 4421 473
rect 4387 371 4421 405
rect 4845 1595 4879 1629
rect 4845 1527 4879 1557
rect 4845 1523 4879 1527
rect 4845 1459 4879 1485
rect 4845 1451 4879 1459
rect 4845 1391 4879 1413
rect 4845 1379 4879 1391
rect 4845 1323 4879 1341
rect 4845 1307 4879 1323
rect 4845 1255 4879 1269
rect 4845 1235 4879 1255
rect 4845 1187 4879 1197
rect 4845 1163 4879 1187
rect 4845 1119 4879 1125
rect 4845 1091 4879 1119
rect 4845 1051 4879 1053
rect 4845 1019 4879 1051
rect 4845 949 4879 981
rect 4845 947 4879 949
rect 4845 881 4879 909
rect 4845 875 4879 881
rect 4845 813 4879 837
rect 4845 803 4879 813
rect 4845 745 4879 765
rect 4845 731 4879 745
rect 4845 677 4879 693
rect 4845 659 4879 677
rect 4845 609 4879 621
rect 4845 587 4879 609
rect 4845 541 4879 549
rect 4845 515 4879 541
rect 4845 473 4879 477
rect 4845 443 4879 473
rect 4845 371 4879 405
rect 5303 1595 5337 1629
rect 5303 1527 5337 1557
rect 5303 1523 5337 1527
rect 5303 1459 5337 1485
rect 5303 1451 5337 1459
rect 5303 1391 5337 1413
rect 5303 1379 5337 1391
rect 5303 1323 5337 1341
rect 5303 1307 5337 1323
rect 5303 1255 5337 1269
rect 5303 1235 5337 1255
rect 5303 1187 5337 1197
rect 5303 1163 5337 1187
rect 5303 1119 5337 1125
rect 5303 1091 5337 1119
rect 5303 1051 5337 1053
rect 5303 1019 5337 1051
rect 5303 949 5337 981
rect 5303 947 5337 949
rect 5303 881 5337 909
rect 5303 875 5337 881
rect 5303 813 5337 837
rect 5303 803 5337 813
rect 5303 745 5337 765
rect 5303 731 5337 745
rect 5303 677 5337 693
rect 5303 659 5337 677
rect 5303 609 5337 621
rect 5303 587 5337 609
rect 5303 541 5337 549
rect 5303 515 5337 541
rect 5303 473 5337 477
rect 5303 443 5337 473
rect 5303 371 5337 405
rect 5761 1595 5795 1629
rect 5761 1527 5795 1557
rect 5761 1523 5795 1527
rect 5761 1459 5795 1485
rect 5761 1451 5795 1459
rect 5761 1391 5795 1413
rect 5761 1379 5795 1391
rect 5761 1323 5795 1341
rect 5761 1307 5795 1323
rect 5761 1255 5795 1269
rect 5761 1235 5795 1255
rect 5761 1187 5795 1197
rect 5761 1163 5795 1187
rect 5761 1119 5795 1125
rect 5761 1091 5795 1119
rect 5761 1051 5795 1053
rect 5761 1019 5795 1051
rect 5761 949 5795 981
rect 5761 947 5795 949
rect 5761 881 5795 909
rect 5761 875 5795 881
rect 5761 813 5795 837
rect 5761 803 5795 813
rect 5761 745 5795 765
rect 5761 731 5795 745
rect 5761 677 5795 693
rect 5761 659 5795 677
rect 5761 609 5795 621
rect 5761 587 5795 609
rect 5761 541 5795 549
rect 5761 515 5795 541
rect 5761 473 5795 477
rect 5761 443 5795 473
rect 5761 371 5795 405
rect 401 -17 435 17
rect 801 -17 835 17
rect 1201 -17 1235 17
rect 1601 -17 1635 17
rect 2001 -17 2035 17
rect 2401 -17 2435 17
rect 2801 -17 2835 17
rect 3201 -17 3235 17
rect 3601 -17 3635 17
rect 4001 -17 4035 17
rect 4401 -17 4435 17
rect 4801 -17 4835 17
rect 5201 -17 5235 17
rect 5601 -17 5635 17
<< metal1 >>
rect 120 1897 5842 1940
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3201 1897
rect 3235 1863 3601 1897
rect 3635 1863 4001 1897
rect 4035 1863 4401 1897
rect 4435 1863 4801 1897
rect 4835 1863 5201 1897
rect 5235 1863 5601 1897
rect 5635 1863 5842 1897
rect 120 1820 5842 1863
rect 259 1629 305 1645
rect 259 1595 265 1629
rect 299 1595 305 1629
rect 259 1557 305 1595
rect 259 1523 265 1557
rect 299 1523 305 1557
rect 259 1485 305 1523
rect 259 1451 265 1485
rect 299 1451 305 1485
rect 259 1413 305 1451
rect 259 1379 265 1413
rect 299 1379 305 1413
rect 259 1341 305 1379
rect 259 1307 265 1341
rect 299 1307 305 1341
rect 259 1269 305 1307
rect 259 1235 265 1269
rect 299 1235 305 1269
rect 259 1197 305 1235
rect 259 1163 265 1197
rect 299 1163 305 1197
rect 259 1125 305 1163
rect 259 1091 265 1125
rect 299 1091 305 1125
rect 259 1053 305 1091
rect 259 1019 265 1053
rect 299 1019 305 1053
rect 259 981 305 1019
rect 259 947 265 981
rect 299 947 305 981
rect 259 909 305 947
rect 259 875 265 909
rect 299 875 305 909
rect 259 837 305 875
rect 259 803 265 837
rect 299 803 305 837
rect 259 765 305 803
rect 259 731 265 765
rect 299 731 305 765
rect 259 693 305 731
rect 259 659 265 693
rect 299 659 305 693
rect 259 621 305 659
rect 259 587 265 621
rect 299 587 305 621
rect 259 549 305 587
rect 259 515 265 549
rect 299 515 305 549
rect 259 477 305 515
rect 259 443 265 477
rect 299 443 305 477
rect 259 405 305 443
rect 259 371 265 405
rect 299 371 305 405
rect 259 355 305 371
rect 717 1629 763 1645
rect 717 1595 723 1629
rect 757 1595 763 1629
rect 717 1557 763 1595
rect 717 1523 723 1557
rect 757 1523 763 1557
rect 717 1485 763 1523
rect 717 1451 723 1485
rect 757 1451 763 1485
rect 717 1413 763 1451
rect 717 1379 723 1413
rect 757 1379 763 1413
rect 717 1341 763 1379
rect 717 1307 723 1341
rect 757 1307 763 1341
rect 717 1269 763 1307
rect 717 1235 723 1269
rect 757 1235 763 1269
rect 717 1197 763 1235
rect 717 1163 723 1197
rect 757 1163 763 1197
rect 717 1125 763 1163
rect 717 1091 723 1125
rect 757 1091 763 1125
rect 717 1053 763 1091
rect 717 1019 723 1053
rect 757 1019 763 1053
rect 717 981 763 1019
rect 717 947 723 981
rect 757 947 763 981
rect 717 909 763 947
rect 717 875 723 909
rect 757 875 763 909
rect 717 837 763 875
rect 717 803 723 837
rect 757 803 763 837
rect 717 765 763 803
rect 717 731 723 765
rect 757 731 763 765
rect 717 693 763 731
rect 717 659 723 693
rect 757 659 763 693
rect 717 621 763 659
rect 717 587 723 621
rect 757 587 763 621
rect 717 549 763 587
rect 717 515 723 549
rect 757 515 763 549
rect 717 477 763 515
rect 717 443 723 477
rect 757 443 763 477
rect 717 405 763 443
rect 717 371 723 405
rect 757 371 763 405
rect 717 355 763 371
rect 1175 1629 1221 1645
rect 1175 1595 1181 1629
rect 1215 1595 1221 1629
rect 1175 1557 1221 1595
rect 1175 1523 1181 1557
rect 1215 1523 1221 1557
rect 1175 1485 1221 1523
rect 1175 1451 1181 1485
rect 1215 1451 1221 1485
rect 1175 1413 1221 1451
rect 1175 1379 1181 1413
rect 1215 1379 1221 1413
rect 1175 1341 1221 1379
rect 1175 1307 1181 1341
rect 1215 1307 1221 1341
rect 1175 1269 1221 1307
rect 1175 1235 1181 1269
rect 1215 1235 1221 1269
rect 1175 1197 1221 1235
rect 1175 1163 1181 1197
rect 1215 1163 1221 1197
rect 1175 1125 1221 1163
rect 1175 1091 1181 1125
rect 1215 1091 1221 1125
rect 1175 1053 1221 1091
rect 1175 1019 1181 1053
rect 1215 1019 1221 1053
rect 1175 981 1221 1019
rect 1175 947 1181 981
rect 1215 947 1221 981
rect 1175 909 1221 947
rect 1175 875 1181 909
rect 1215 875 1221 909
rect 1175 837 1221 875
rect 1175 803 1181 837
rect 1215 803 1221 837
rect 1175 765 1221 803
rect 1175 731 1181 765
rect 1215 731 1221 765
rect 1175 693 1221 731
rect 1175 659 1181 693
rect 1215 659 1221 693
rect 1175 621 1221 659
rect 1175 587 1181 621
rect 1215 587 1221 621
rect 1175 549 1221 587
rect 1175 515 1181 549
rect 1215 515 1221 549
rect 1175 477 1221 515
rect 1175 443 1181 477
rect 1215 443 1221 477
rect 1175 405 1221 443
rect 1175 371 1181 405
rect 1215 371 1221 405
rect 1175 355 1221 371
rect 1633 1629 1679 1645
rect 1633 1595 1639 1629
rect 1673 1595 1679 1629
rect 1633 1557 1679 1595
rect 1633 1523 1639 1557
rect 1673 1523 1679 1557
rect 1633 1485 1679 1523
rect 1633 1451 1639 1485
rect 1673 1451 1679 1485
rect 1633 1413 1679 1451
rect 1633 1379 1639 1413
rect 1673 1379 1679 1413
rect 1633 1341 1679 1379
rect 1633 1307 1639 1341
rect 1673 1307 1679 1341
rect 1633 1269 1679 1307
rect 1633 1235 1639 1269
rect 1673 1235 1679 1269
rect 1633 1197 1679 1235
rect 1633 1163 1639 1197
rect 1673 1163 1679 1197
rect 1633 1125 1679 1163
rect 1633 1091 1639 1125
rect 1673 1091 1679 1125
rect 1633 1053 1679 1091
rect 1633 1019 1639 1053
rect 1673 1019 1679 1053
rect 1633 981 1679 1019
rect 1633 947 1639 981
rect 1673 947 1679 981
rect 1633 909 1679 947
rect 1633 875 1639 909
rect 1673 875 1679 909
rect 1633 837 1679 875
rect 1633 803 1639 837
rect 1673 803 1679 837
rect 1633 765 1679 803
rect 1633 731 1639 765
rect 1673 731 1679 765
rect 1633 693 1679 731
rect 1633 659 1639 693
rect 1673 659 1679 693
rect 1633 621 1679 659
rect 1633 587 1639 621
rect 1673 587 1679 621
rect 1633 549 1679 587
rect 1633 515 1639 549
rect 1673 515 1679 549
rect 1633 477 1679 515
rect 1633 443 1639 477
rect 1673 443 1679 477
rect 1633 405 1679 443
rect 1633 371 1639 405
rect 1673 371 1679 405
rect 1633 355 1679 371
rect 2091 1629 2137 1645
rect 2091 1595 2097 1629
rect 2131 1595 2137 1629
rect 2091 1557 2137 1595
rect 2091 1523 2097 1557
rect 2131 1523 2137 1557
rect 2091 1485 2137 1523
rect 2091 1451 2097 1485
rect 2131 1451 2137 1485
rect 2091 1413 2137 1451
rect 2091 1379 2097 1413
rect 2131 1379 2137 1413
rect 2091 1341 2137 1379
rect 2091 1307 2097 1341
rect 2131 1307 2137 1341
rect 2091 1269 2137 1307
rect 2091 1235 2097 1269
rect 2131 1235 2137 1269
rect 2091 1197 2137 1235
rect 2091 1163 2097 1197
rect 2131 1163 2137 1197
rect 2091 1125 2137 1163
rect 2091 1091 2097 1125
rect 2131 1091 2137 1125
rect 2091 1053 2137 1091
rect 2091 1019 2097 1053
rect 2131 1019 2137 1053
rect 2091 981 2137 1019
rect 2091 947 2097 981
rect 2131 947 2137 981
rect 2091 909 2137 947
rect 2091 875 2097 909
rect 2131 875 2137 909
rect 2091 837 2137 875
rect 2091 803 2097 837
rect 2131 803 2137 837
rect 2091 765 2137 803
rect 2091 731 2097 765
rect 2131 731 2137 765
rect 2091 693 2137 731
rect 2091 659 2097 693
rect 2131 659 2137 693
rect 2091 621 2137 659
rect 2091 587 2097 621
rect 2131 587 2137 621
rect 2091 549 2137 587
rect 2091 515 2097 549
rect 2131 515 2137 549
rect 2091 477 2137 515
rect 2091 443 2097 477
rect 2131 443 2137 477
rect 2091 405 2137 443
rect 2091 371 2097 405
rect 2131 371 2137 405
rect 2091 355 2137 371
rect 2549 1629 2595 1645
rect 2549 1595 2555 1629
rect 2589 1595 2595 1629
rect 2549 1557 2595 1595
rect 2549 1523 2555 1557
rect 2589 1523 2595 1557
rect 2549 1485 2595 1523
rect 2549 1451 2555 1485
rect 2589 1451 2595 1485
rect 2549 1413 2595 1451
rect 2549 1379 2555 1413
rect 2589 1379 2595 1413
rect 2549 1341 2595 1379
rect 2549 1307 2555 1341
rect 2589 1307 2595 1341
rect 2549 1269 2595 1307
rect 2549 1235 2555 1269
rect 2589 1235 2595 1269
rect 2549 1197 2595 1235
rect 2549 1163 2555 1197
rect 2589 1163 2595 1197
rect 2549 1125 2595 1163
rect 2549 1091 2555 1125
rect 2589 1091 2595 1125
rect 2549 1053 2595 1091
rect 2549 1019 2555 1053
rect 2589 1019 2595 1053
rect 2549 981 2595 1019
rect 2549 947 2555 981
rect 2589 947 2595 981
rect 2549 909 2595 947
rect 2549 875 2555 909
rect 2589 875 2595 909
rect 2549 837 2595 875
rect 2549 803 2555 837
rect 2589 803 2595 837
rect 2549 765 2595 803
rect 2549 731 2555 765
rect 2589 731 2595 765
rect 2549 693 2595 731
rect 2549 659 2555 693
rect 2589 659 2595 693
rect 2549 621 2595 659
rect 2549 587 2555 621
rect 2589 587 2595 621
rect 2549 549 2595 587
rect 2549 515 2555 549
rect 2589 515 2595 549
rect 2549 477 2595 515
rect 2549 443 2555 477
rect 2589 443 2595 477
rect 2549 405 2595 443
rect 2549 371 2555 405
rect 2589 371 2595 405
rect 2549 355 2595 371
rect 3007 1629 3053 1645
rect 3007 1595 3013 1629
rect 3047 1595 3053 1629
rect 3007 1557 3053 1595
rect 3007 1523 3013 1557
rect 3047 1523 3053 1557
rect 3007 1485 3053 1523
rect 3007 1451 3013 1485
rect 3047 1451 3053 1485
rect 3007 1413 3053 1451
rect 3007 1379 3013 1413
rect 3047 1379 3053 1413
rect 3007 1341 3053 1379
rect 3007 1307 3013 1341
rect 3047 1307 3053 1341
rect 3007 1269 3053 1307
rect 3007 1235 3013 1269
rect 3047 1235 3053 1269
rect 3007 1197 3053 1235
rect 3007 1163 3013 1197
rect 3047 1163 3053 1197
rect 3007 1125 3053 1163
rect 3007 1091 3013 1125
rect 3047 1091 3053 1125
rect 3007 1053 3053 1091
rect 3007 1019 3013 1053
rect 3047 1019 3053 1053
rect 3007 981 3053 1019
rect 3007 947 3013 981
rect 3047 947 3053 981
rect 3007 909 3053 947
rect 3007 875 3013 909
rect 3047 875 3053 909
rect 3007 837 3053 875
rect 3007 803 3013 837
rect 3047 803 3053 837
rect 3007 765 3053 803
rect 3007 731 3013 765
rect 3047 731 3053 765
rect 3007 693 3053 731
rect 3007 659 3013 693
rect 3047 659 3053 693
rect 3007 621 3053 659
rect 3007 587 3013 621
rect 3047 587 3053 621
rect 3007 549 3053 587
rect 3007 515 3013 549
rect 3047 515 3053 549
rect 3007 477 3053 515
rect 3007 443 3013 477
rect 3047 443 3053 477
rect 3007 405 3053 443
rect 3007 371 3013 405
rect 3047 371 3053 405
rect 3007 355 3053 371
rect 3465 1629 3511 1645
rect 3465 1595 3471 1629
rect 3505 1595 3511 1629
rect 3465 1557 3511 1595
rect 3465 1523 3471 1557
rect 3505 1523 3511 1557
rect 3465 1485 3511 1523
rect 3465 1451 3471 1485
rect 3505 1451 3511 1485
rect 3465 1413 3511 1451
rect 3465 1379 3471 1413
rect 3505 1379 3511 1413
rect 3465 1341 3511 1379
rect 3465 1307 3471 1341
rect 3505 1307 3511 1341
rect 3465 1269 3511 1307
rect 3465 1235 3471 1269
rect 3505 1235 3511 1269
rect 3465 1197 3511 1235
rect 3465 1163 3471 1197
rect 3505 1163 3511 1197
rect 3465 1125 3511 1163
rect 3465 1091 3471 1125
rect 3505 1091 3511 1125
rect 3465 1053 3511 1091
rect 3465 1019 3471 1053
rect 3505 1019 3511 1053
rect 3465 981 3511 1019
rect 3465 947 3471 981
rect 3505 947 3511 981
rect 3465 909 3511 947
rect 3465 875 3471 909
rect 3505 875 3511 909
rect 3465 837 3511 875
rect 3465 803 3471 837
rect 3505 803 3511 837
rect 3465 765 3511 803
rect 3465 731 3471 765
rect 3505 731 3511 765
rect 3465 693 3511 731
rect 3465 659 3471 693
rect 3505 659 3511 693
rect 3465 621 3511 659
rect 3465 587 3471 621
rect 3505 587 3511 621
rect 3465 549 3511 587
rect 3465 515 3471 549
rect 3505 515 3511 549
rect 3465 477 3511 515
rect 3465 443 3471 477
rect 3505 443 3511 477
rect 3465 405 3511 443
rect 3465 371 3471 405
rect 3505 371 3511 405
rect 3465 355 3511 371
rect 3923 1629 3969 1645
rect 3923 1595 3929 1629
rect 3963 1595 3969 1629
rect 3923 1557 3969 1595
rect 3923 1523 3929 1557
rect 3963 1523 3969 1557
rect 3923 1485 3969 1523
rect 3923 1451 3929 1485
rect 3963 1451 3969 1485
rect 3923 1413 3969 1451
rect 3923 1379 3929 1413
rect 3963 1379 3969 1413
rect 3923 1341 3969 1379
rect 3923 1307 3929 1341
rect 3963 1307 3969 1341
rect 3923 1269 3969 1307
rect 3923 1235 3929 1269
rect 3963 1235 3969 1269
rect 3923 1197 3969 1235
rect 3923 1163 3929 1197
rect 3963 1163 3969 1197
rect 3923 1125 3969 1163
rect 3923 1091 3929 1125
rect 3963 1091 3969 1125
rect 3923 1053 3969 1091
rect 3923 1019 3929 1053
rect 3963 1019 3969 1053
rect 3923 981 3969 1019
rect 3923 947 3929 981
rect 3963 947 3969 981
rect 3923 909 3969 947
rect 3923 875 3929 909
rect 3963 875 3969 909
rect 3923 837 3969 875
rect 3923 803 3929 837
rect 3963 803 3969 837
rect 3923 765 3969 803
rect 3923 731 3929 765
rect 3963 731 3969 765
rect 3923 693 3969 731
rect 3923 659 3929 693
rect 3963 659 3969 693
rect 3923 621 3969 659
rect 3923 587 3929 621
rect 3963 587 3969 621
rect 3923 549 3969 587
rect 3923 515 3929 549
rect 3963 515 3969 549
rect 3923 477 3969 515
rect 3923 443 3929 477
rect 3963 443 3969 477
rect 3923 405 3969 443
rect 3923 371 3929 405
rect 3963 371 3969 405
rect 3923 355 3969 371
rect 4381 1629 4427 1645
rect 4381 1595 4387 1629
rect 4421 1595 4427 1629
rect 4381 1557 4427 1595
rect 4381 1523 4387 1557
rect 4421 1523 4427 1557
rect 4381 1485 4427 1523
rect 4381 1451 4387 1485
rect 4421 1451 4427 1485
rect 4381 1413 4427 1451
rect 4381 1379 4387 1413
rect 4421 1379 4427 1413
rect 4381 1341 4427 1379
rect 4381 1307 4387 1341
rect 4421 1307 4427 1341
rect 4381 1269 4427 1307
rect 4381 1235 4387 1269
rect 4421 1235 4427 1269
rect 4381 1197 4427 1235
rect 4381 1163 4387 1197
rect 4421 1163 4427 1197
rect 4381 1125 4427 1163
rect 4381 1091 4387 1125
rect 4421 1091 4427 1125
rect 4381 1053 4427 1091
rect 4381 1019 4387 1053
rect 4421 1019 4427 1053
rect 4381 981 4427 1019
rect 4381 947 4387 981
rect 4421 947 4427 981
rect 4381 909 4427 947
rect 4381 875 4387 909
rect 4421 875 4427 909
rect 4381 837 4427 875
rect 4381 803 4387 837
rect 4421 803 4427 837
rect 4381 765 4427 803
rect 4381 731 4387 765
rect 4421 731 4427 765
rect 4381 693 4427 731
rect 4381 659 4387 693
rect 4421 659 4427 693
rect 4381 621 4427 659
rect 4381 587 4387 621
rect 4421 587 4427 621
rect 4381 549 4427 587
rect 4381 515 4387 549
rect 4421 515 4427 549
rect 4381 477 4427 515
rect 4381 443 4387 477
rect 4421 443 4427 477
rect 4381 405 4427 443
rect 4381 371 4387 405
rect 4421 371 4427 405
rect 4381 355 4427 371
rect 4839 1629 4885 1645
rect 4839 1595 4845 1629
rect 4879 1595 4885 1629
rect 4839 1557 4885 1595
rect 4839 1523 4845 1557
rect 4879 1523 4885 1557
rect 4839 1485 4885 1523
rect 4839 1451 4845 1485
rect 4879 1451 4885 1485
rect 4839 1413 4885 1451
rect 4839 1379 4845 1413
rect 4879 1379 4885 1413
rect 4839 1341 4885 1379
rect 4839 1307 4845 1341
rect 4879 1307 4885 1341
rect 4839 1269 4885 1307
rect 4839 1235 4845 1269
rect 4879 1235 4885 1269
rect 4839 1197 4885 1235
rect 4839 1163 4845 1197
rect 4879 1163 4885 1197
rect 4839 1125 4885 1163
rect 4839 1091 4845 1125
rect 4879 1091 4885 1125
rect 4839 1053 4885 1091
rect 4839 1019 4845 1053
rect 4879 1019 4885 1053
rect 4839 981 4885 1019
rect 4839 947 4845 981
rect 4879 947 4885 981
rect 4839 909 4885 947
rect 4839 875 4845 909
rect 4879 875 4885 909
rect 4839 837 4885 875
rect 4839 803 4845 837
rect 4879 803 4885 837
rect 4839 765 4885 803
rect 4839 731 4845 765
rect 4879 731 4885 765
rect 4839 693 4885 731
rect 4839 659 4845 693
rect 4879 659 4885 693
rect 4839 621 4885 659
rect 4839 587 4845 621
rect 4879 587 4885 621
rect 4839 549 4885 587
rect 4839 515 4845 549
rect 4879 515 4885 549
rect 4839 477 4885 515
rect 4839 443 4845 477
rect 4879 443 4885 477
rect 4839 405 4885 443
rect 4839 371 4845 405
rect 4879 371 4885 405
rect 4839 355 4885 371
rect 5297 1629 5343 1645
rect 5297 1595 5303 1629
rect 5337 1595 5343 1629
rect 5297 1557 5343 1595
rect 5297 1523 5303 1557
rect 5337 1523 5343 1557
rect 5297 1485 5343 1523
rect 5297 1451 5303 1485
rect 5337 1451 5343 1485
rect 5297 1413 5343 1451
rect 5297 1379 5303 1413
rect 5337 1379 5343 1413
rect 5297 1341 5343 1379
rect 5297 1307 5303 1341
rect 5337 1307 5343 1341
rect 5297 1269 5343 1307
rect 5297 1235 5303 1269
rect 5337 1235 5343 1269
rect 5297 1197 5343 1235
rect 5297 1163 5303 1197
rect 5337 1163 5343 1197
rect 5297 1125 5343 1163
rect 5297 1091 5303 1125
rect 5337 1091 5343 1125
rect 5297 1053 5343 1091
rect 5297 1019 5303 1053
rect 5337 1019 5343 1053
rect 5297 981 5343 1019
rect 5297 947 5303 981
rect 5337 947 5343 981
rect 5297 909 5343 947
rect 5297 875 5303 909
rect 5337 875 5343 909
rect 5297 837 5343 875
rect 5297 803 5303 837
rect 5337 803 5343 837
rect 5297 765 5343 803
rect 5297 731 5303 765
rect 5337 731 5343 765
rect 5297 693 5343 731
rect 5297 659 5303 693
rect 5337 659 5343 693
rect 5297 621 5343 659
rect 5297 587 5303 621
rect 5337 587 5343 621
rect 5297 549 5343 587
rect 5297 515 5303 549
rect 5337 515 5343 549
rect 5297 477 5343 515
rect 5297 443 5303 477
rect 5337 443 5343 477
rect 5297 405 5343 443
rect 5297 371 5303 405
rect 5337 371 5343 405
rect 5297 355 5343 371
rect 5755 1629 5801 1645
rect 5755 1595 5761 1629
rect 5795 1595 5801 1629
rect 5755 1557 5801 1595
rect 5755 1523 5761 1557
rect 5795 1523 5801 1557
rect 5755 1485 5801 1523
rect 5755 1451 5761 1485
rect 5795 1451 5801 1485
rect 5755 1413 5801 1451
rect 5755 1379 5761 1413
rect 5795 1379 5801 1413
rect 5755 1341 5801 1379
rect 5755 1307 5761 1341
rect 5795 1307 5801 1341
rect 5755 1269 5801 1307
rect 5755 1235 5761 1269
rect 5795 1235 5801 1269
rect 5755 1197 5801 1235
rect 5755 1163 5761 1197
rect 5795 1163 5801 1197
rect 5755 1125 5801 1163
rect 5755 1091 5761 1125
rect 5795 1091 5801 1125
rect 5755 1053 5801 1091
rect 5755 1019 5761 1053
rect 5795 1019 5801 1053
rect 5755 981 5801 1019
rect 5755 947 5761 981
rect 5795 947 5801 981
rect 5755 909 5801 947
rect 5755 875 5761 909
rect 5795 875 5801 909
rect 5755 837 5801 875
rect 5755 803 5761 837
rect 5795 803 5801 837
rect 5755 765 5801 803
rect 5755 731 5761 765
rect 5795 731 5801 765
rect 5755 693 5801 731
rect 5755 659 5761 693
rect 5795 659 5801 693
rect 5755 621 5801 659
rect 5755 587 5761 621
rect 5795 587 5801 621
rect 5755 549 5801 587
rect 5755 515 5761 549
rect 5795 515 5801 549
rect 5755 477 5801 515
rect 5755 443 5761 477
rect 5795 443 5801 477
rect 5755 405 5801 443
rect 5755 371 5761 405
rect 5795 371 5801 405
rect 5755 355 5801 371
rect 120 17 5842 60
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3201 17
rect 3235 -17 3601 17
rect 3635 -17 4001 17
rect 4035 -17 4401 17
rect 4435 -17 4801 17
rect 4835 -17 5201 17
rect 5235 -17 5601 17
rect 5635 -17 5842 17
rect 120 -60 5842 -17
<< labels >>
flabel locali s 5782 104 5842 164 1 FreeSans 1952 0 0 0 GATE
port 1 nsew
flabel locali s 5782 1690 5842 1730 1 FreeSans 1952 0 0 0 SOURCE
port 2 nsew
flabel locali s 5782 210 5842 270 1 FreeSans 1952 0 0 0 DRAIN
port 3 nsew
flabel nwell s 120 1850 180 1910 1 FreeSans 1952 0 0 0 VPWR
port 4 nsew
flabel metal1 s 120 -30 278 30 1 FreeSans 1952 0 0 0 VGND
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 5963 1880
<< end >>
