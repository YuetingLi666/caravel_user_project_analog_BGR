magic
tech sky130A
timestamp 1655816534
<< metal1 >>
rect -13 13 13 16
rect -13 -16 13 -13
<< via1 >>
rect -13 -13 13 13
<< metal2 >>
rect -13 13 13 16
rect -13 -16 13 -13
<< end >>
