magic
tech sky130A
magscale 1 2
timestamp 1654901230
<< pwell >>
rect 120 1457 1460 1610
rect 120 423 273 1457
rect 1307 423 1460 1457
rect 120 270 1460 423
<< nbase >>
rect 273 423 1307 1457
<< pdiff >>
rect 450 1228 1130 1280
rect 450 1194 504 1228
rect 538 1194 594 1228
rect 628 1194 684 1228
rect 718 1194 774 1228
rect 808 1194 864 1228
rect 898 1194 954 1228
rect 988 1194 1044 1228
rect 1078 1194 1130 1228
rect 450 1138 1130 1194
rect 450 1104 504 1138
rect 538 1104 594 1138
rect 628 1104 684 1138
rect 718 1104 774 1138
rect 808 1104 864 1138
rect 898 1104 954 1138
rect 988 1104 1044 1138
rect 1078 1104 1130 1138
rect 450 1048 1130 1104
rect 450 1014 504 1048
rect 538 1014 594 1048
rect 628 1014 684 1048
rect 718 1014 774 1048
rect 808 1014 864 1048
rect 898 1014 954 1048
rect 988 1014 1044 1048
rect 1078 1014 1130 1048
rect 450 958 1130 1014
rect 450 924 504 958
rect 538 924 594 958
rect 628 924 684 958
rect 718 924 774 958
rect 808 924 864 958
rect 898 924 954 958
rect 988 924 1044 958
rect 1078 924 1130 958
rect 450 868 1130 924
rect 450 834 504 868
rect 538 834 594 868
rect 628 834 684 868
rect 718 834 774 868
rect 808 834 864 868
rect 898 834 954 868
rect 988 834 1044 868
rect 1078 834 1130 868
rect 450 778 1130 834
rect 450 744 504 778
rect 538 744 594 778
rect 628 744 684 778
rect 718 744 774 778
rect 808 744 864 778
rect 898 744 954 778
rect 988 744 1044 778
rect 1078 744 1130 778
rect 450 688 1130 744
rect 450 654 504 688
rect 538 654 594 688
rect 628 654 684 688
rect 718 654 774 688
rect 808 654 864 688
rect 898 654 954 688
rect 988 654 1044 688
rect 1078 654 1130 688
rect 450 600 1130 654
<< pdiffc >>
rect 504 1194 538 1228
rect 594 1194 628 1228
rect 684 1194 718 1228
rect 774 1194 808 1228
rect 864 1194 898 1228
rect 954 1194 988 1228
rect 1044 1194 1078 1228
rect 504 1104 538 1138
rect 594 1104 628 1138
rect 684 1104 718 1138
rect 774 1104 808 1138
rect 864 1104 898 1138
rect 954 1104 988 1138
rect 1044 1104 1078 1138
rect 504 1014 538 1048
rect 594 1014 628 1048
rect 684 1014 718 1048
rect 774 1014 808 1048
rect 864 1014 898 1048
rect 954 1014 988 1048
rect 1044 1014 1078 1048
rect 504 924 538 958
rect 594 924 628 958
rect 684 924 718 958
rect 774 924 808 958
rect 864 924 898 958
rect 954 924 988 958
rect 1044 924 1078 958
rect 504 834 538 868
rect 594 834 628 868
rect 684 834 718 868
rect 774 834 808 868
rect 864 834 898 868
rect 954 834 988 868
rect 1044 834 1078 868
rect 504 744 538 778
rect 594 744 628 778
rect 684 744 718 778
rect 774 744 808 778
rect 864 744 898 778
rect 954 744 988 778
rect 1044 744 1078 778
rect 504 654 538 688
rect 594 654 628 688
rect 684 654 718 688
rect 774 654 808 688
rect 864 654 898 688
rect 954 654 988 688
rect 1044 654 1078 688
<< psubdiff >>
rect 146 1549 1434 1584
rect 146 1526 276 1549
rect 146 1492 180 1526
rect 214 1515 276 1526
rect 310 1515 366 1549
rect 400 1515 456 1549
rect 490 1515 546 1549
rect 580 1515 636 1549
rect 670 1515 726 1549
rect 760 1515 816 1549
rect 850 1515 906 1549
rect 940 1515 996 1549
rect 1030 1515 1086 1549
rect 1120 1515 1176 1549
rect 1210 1515 1266 1549
rect 1300 1526 1434 1549
rect 1300 1515 1367 1526
rect 214 1492 1367 1515
rect 1401 1492 1434 1526
rect 146 1483 1434 1492
rect 146 1436 247 1483
rect 146 1402 180 1436
rect 214 1402 247 1436
rect 1333 1436 1434 1483
rect 146 1346 247 1402
rect 146 1312 180 1346
rect 214 1312 247 1346
rect 146 1256 247 1312
rect 146 1222 180 1256
rect 214 1222 247 1256
rect 146 1166 247 1222
rect 146 1132 180 1166
rect 214 1132 247 1166
rect 146 1076 247 1132
rect 146 1042 180 1076
rect 214 1042 247 1076
rect 146 986 247 1042
rect 146 952 180 986
rect 214 952 247 986
rect 146 896 247 952
rect 146 862 180 896
rect 214 862 247 896
rect 146 806 247 862
rect 146 772 180 806
rect 214 772 247 806
rect 146 716 247 772
rect 146 682 180 716
rect 214 682 247 716
rect 146 626 247 682
rect 146 592 180 626
rect 214 592 247 626
rect 146 536 247 592
rect 146 502 180 536
rect 214 502 247 536
rect 146 446 247 502
rect 1333 1402 1367 1436
rect 1401 1402 1434 1436
rect 1333 1346 1434 1402
rect 1333 1312 1367 1346
rect 1401 1312 1434 1346
rect 1333 1256 1434 1312
rect 1333 1222 1367 1256
rect 1401 1222 1434 1256
rect 1333 1166 1434 1222
rect 1333 1132 1367 1166
rect 1401 1132 1434 1166
rect 1333 1076 1434 1132
rect 1333 1042 1367 1076
rect 1401 1042 1434 1076
rect 1333 986 1434 1042
rect 1333 952 1367 986
rect 1401 952 1434 986
rect 1333 896 1434 952
rect 1333 862 1367 896
rect 1401 862 1434 896
rect 1333 806 1434 862
rect 1333 772 1367 806
rect 1401 772 1434 806
rect 1333 716 1434 772
rect 1333 682 1367 716
rect 1401 682 1434 716
rect 1333 626 1434 682
rect 1333 592 1367 626
rect 1401 592 1434 626
rect 1333 536 1434 592
rect 1333 502 1367 536
rect 1401 502 1434 536
rect 146 412 180 446
rect 214 412 247 446
rect 146 397 247 412
rect 1333 446 1434 502
rect 1333 412 1367 446
rect 1401 412 1434 446
rect 1333 397 1434 412
rect 146 362 1434 397
rect 146 328 276 362
rect 310 328 366 362
rect 400 328 456 362
rect 490 328 546 362
rect 580 328 636 362
rect 670 328 726 362
rect 760 328 816 362
rect 850 328 906 362
rect 940 328 996 362
rect 1030 328 1086 362
rect 1120 328 1176 362
rect 1210 328 1266 362
rect 1300 328 1434 362
rect 146 296 1434 328
<< nsubdiff >>
rect 309 1402 1271 1421
rect 309 1368 440 1402
rect 474 1368 530 1402
rect 564 1368 620 1402
rect 654 1368 710 1402
rect 744 1368 800 1402
rect 834 1368 890 1402
rect 924 1368 980 1402
rect 1014 1368 1070 1402
rect 1104 1368 1160 1402
rect 1194 1368 1271 1402
rect 309 1349 1271 1368
rect 309 1345 381 1349
rect 309 1311 328 1345
rect 362 1311 381 1345
rect 309 1255 381 1311
rect 1199 1326 1271 1349
rect 1199 1292 1218 1326
rect 1252 1292 1271 1326
rect 309 1221 328 1255
rect 362 1221 381 1255
rect 309 1165 381 1221
rect 309 1131 328 1165
rect 362 1131 381 1165
rect 309 1075 381 1131
rect 309 1041 328 1075
rect 362 1041 381 1075
rect 309 985 381 1041
rect 309 951 328 985
rect 362 951 381 985
rect 309 895 381 951
rect 309 861 328 895
rect 362 861 381 895
rect 309 805 381 861
rect 309 771 328 805
rect 362 771 381 805
rect 309 715 381 771
rect 309 681 328 715
rect 362 681 381 715
rect 309 625 381 681
rect 309 591 328 625
rect 362 591 381 625
rect 1199 1236 1271 1292
rect 1199 1202 1218 1236
rect 1252 1202 1271 1236
rect 1199 1146 1271 1202
rect 1199 1112 1218 1146
rect 1252 1112 1271 1146
rect 1199 1056 1271 1112
rect 1199 1022 1218 1056
rect 1252 1022 1271 1056
rect 1199 966 1271 1022
rect 1199 932 1218 966
rect 1252 932 1271 966
rect 1199 876 1271 932
rect 1199 842 1218 876
rect 1252 842 1271 876
rect 1199 786 1271 842
rect 1199 752 1218 786
rect 1252 752 1271 786
rect 1199 696 1271 752
rect 1199 662 1218 696
rect 1252 662 1271 696
rect 1199 606 1271 662
rect 309 531 381 591
rect 1199 572 1218 606
rect 1252 572 1271 606
rect 1199 531 1271 572
rect 309 512 1271 531
rect 309 478 406 512
rect 440 478 496 512
rect 530 478 586 512
rect 620 478 676 512
rect 710 478 766 512
rect 800 478 856 512
rect 890 478 946 512
rect 980 478 1036 512
rect 1070 478 1126 512
rect 1160 478 1271 512
rect 309 459 1271 478
<< psubdiffcont >>
rect 180 1492 214 1526
rect 276 1515 310 1549
rect 366 1515 400 1549
rect 456 1515 490 1549
rect 546 1515 580 1549
rect 636 1515 670 1549
rect 726 1515 760 1549
rect 816 1515 850 1549
rect 906 1515 940 1549
rect 996 1515 1030 1549
rect 1086 1515 1120 1549
rect 1176 1515 1210 1549
rect 1266 1515 1300 1549
rect 1367 1492 1401 1526
rect 180 1402 214 1436
rect 180 1312 214 1346
rect 180 1222 214 1256
rect 180 1132 214 1166
rect 180 1042 214 1076
rect 180 952 214 986
rect 180 862 214 896
rect 180 772 214 806
rect 180 682 214 716
rect 180 592 214 626
rect 180 502 214 536
rect 1367 1402 1401 1436
rect 1367 1312 1401 1346
rect 1367 1222 1401 1256
rect 1367 1132 1401 1166
rect 1367 1042 1401 1076
rect 1367 952 1401 986
rect 1367 862 1401 896
rect 1367 772 1401 806
rect 1367 682 1401 716
rect 1367 592 1401 626
rect 1367 502 1401 536
rect 180 412 214 446
rect 1367 412 1401 446
rect 276 328 310 362
rect 366 328 400 362
rect 456 328 490 362
rect 546 328 580 362
rect 636 328 670 362
rect 726 328 760 362
rect 816 328 850 362
rect 906 328 940 362
rect 996 328 1030 362
rect 1086 328 1120 362
rect 1176 328 1210 362
rect 1266 328 1300 362
<< nsubdiffcont >>
rect 440 1368 474 1402
rect 530 1368 564 1402
rect 620 1368 654 1402
rect 710 1368 744 1402
rect 800 1368 834 1402
rect 890 1368 924 1402
rect 980 1368 1014 1402
rect 1070 1368 1104 1402
rect 1160 1368 1194 1402
rect 328 1311 362 1345
rect 1218 1292 1252 1326
rect 328 1221 362 1255
rect 328 1131 362 1165
rect 328 1041 362 1075
rect 328 951 362 985
rect 328 861 362 895
rect 328 771 362 805
rect 328 681 362 715
rect 328 591 362 625
rect 1218 1202 1252 1236
rect 1218 1112 1252 1146
rect 1218 1022 1252 1056
rect 1218 932 1252 966
rect 1218 842 1252 876
rect 1218 752 1252 786
rect 1218 662 1252 696
rect 1218 572 1252 606
rect 406 478 440 512
rect 496 478 530 512
rect 586 478 620 512
rect 676 478 710 512
rect 766 478 800 512
rect 856 478 890 512
rect 946 478 980 512
rect 1036 478 1070 512
rect 1126 478 1160 512
<< locali >>
rect 120 1897 1460 1910
rect 120 1863 303 1897
rect 337 1863 503 1897
rect 537 1863 703 1897
rect 737 1863 903 1897
rect 937 1863 1103 1897
rect 1137 1863 1303 1897
rect 1337 1863 1460 1897
rect 120 1850 1460 1863
rect 146 1549 1434 1584
rect 146 1526 276 1549
rect 146 1492 180 1526
rect 214 1515 276 1526
rect 310 1515 366 1549
rect 400 1515 456 1549
rect 490 1515 546 1549
rect 580 1515 636 1549
rect 670 1515 726 1549
rect 760 1515 816 1549
rect 850 1515 906 1549
rect 940 1515 996 1549
rect 1030 1515 1086 1549
rect 1120 1515 1176 1549
rect 1210 1515 1266 1549
rect 1300 1526 1434 1549
rect 1300 1515 1367 1526
rect 214 1492 1367 1515
rect 1401 1492 1434 1526
rect 146 1485 1434 1492
rect 146 1436 245 1485
rect 146 1402 180 1436
rect 214 1402 245 1436
rect 1335 1436 1434 1485
rect 146 1346 245 1402
rect 146 1312 180 1346
rect 214 1312 245 1346
rect 146 1256 245 1312
rect 146 1222 180 1256
rect 214 1222 245 1256
rect 146 1166 245 1222
rect 146 1132 180 1166
rect 214 1132 245 1166
rect 146 1076 245 1132
rect 146 1042 180 1076
rect 214 1042 245 1076
rect 146 986 245 1042
rect 146 952 180 986
rect 214 952 245 986
rect 146 896 245 952
rect 146 862 180 896
rect 214 862 245 896
rect 146 806 245 862
rect 146 772 180 806
rect 214 772 245 806
rect 146 716 245 772
rect 146 682 180 716
rect 214 682 245 716
rect 146 626 245 682
rect 146 592 180 626
rect 214 592 245 626
rect 146 536 245 592
rect 146 502 180 536
rect 214 502 245 536
rect 146 446 245 502
rect 309 1402 1271 1421
rect 309 1368 440 1402
rect 474 1368 530 1402
rect 564 1368 620 1402
rect 654 1368 710 1402
rect 744 1368 800 1402
rect 834 1368 890 1402
rect 924 1368 980 1402
rect 1014 1368 1070 1402
rect 1104 1368 1160 1402
rect 1194 1368 1271 1402
rect 309 1349 1271 1368
rect 309 1345 381 1349
rect 309 1311 328 1345
rect 362 1311 381 1345
rect 309 1255 381 1311
rect 1199 1326 1271 1349
rect 1199 1292 1218 1326
rect 1252 1292 1271 1326
rect 309 1221 328 1255
rect 362 1221 381 1255
rect 309 1165 381 1221
rect 309 1131 328 1165
rect 362 1131 381 1165
rect 309 1075 381 1131
rect 309 1041 328 1075
rect 362 1041 381 1075
rect 309 985 381 1041
rect 309 951 328 985
rect 362 951 381 985
rect 309 895 381 951
rect 309 861 328 895
rect 362 861 381 895
rect 309 805 381 861
rect 309 771 328 805
rect 362 771 381 805
rect 309 715 381 771
rect 309 681 328 715
rect 362 681 381 715
rect 309 625 381 681
rect 309 591 328 625
rect 362 591 381 625
rect 443 1228 1137 1287
rect 443 1194 504 1228
rect 538 1200 594 1228
rect 628 1200 684 1228
rect 718 1200 774 1228
rect 550 1194 594 1200
rect 650 1194 684 1200
rect 750 1194 774 1200
rect 808 1200 864 1228
rect 808 1194 816 1200
rect 443 1166 516 1194
rect 550 1166 616 1194
rect 650 1166 716 1194
rect 750 1166 816 1194
rect 850 1194 864 1200
rect 898 1200 954 1228
rect 898 1194 916 1200
rect 850 1166 916 1194
rect 950 1194 954 1200
rect 988 1200 1044 1228
rect 988 1194 1016 1200
rect 1078 1194 1137 1228
rect 950 1166 1016 1194
rect 1050 1166 1137 1194
rect 443 1138 1137 1166
rect 443 1104 504 1138
rect 538 1104 594 1138
rect 628 1104 684 1138
rect 718 1104 774 1138
rect 808 1104 864 1138
rect 898 1104 954 1138
rect 988 1104 1044 1138
rect 1078 1104 1137 1138
rect 443 1100 1137 1104
rect 443 1066 516 1100
rect 550 1066 616 1100
rect 650 1066 716 1100
rect 750 1066 816 1100
rect 850 1066 916 1100
rect 950 1066 1016 1100
rect 1050 1066 1137 1100
rect 443 1048 1137 1066
rect 443 1014 504 1048
rect 538 1014 594 1048
rect 628 1014 684 1048
rect 718 1014 774 1048
rect 808 1014 864 1048
rect 898 1014 954 1048
rect 988 1014 1044 1048
rect 1078 1014 1137 1048
rect 443 1000 1137 1014
rect 443 966 516 1000
rect 550 966 616 1000
rect 650 966 716 1000
rect 750 966 816 1000
rect 850 966 916 1000
rect 950 966 1016 1000
rect 1050 966 1137 1000
rect 443 958 1137 966
rect 443 924 504 958
rect 538 924 594 958
rect 628 924 684 958
rect 718 924 774 958
rect 808 924 864 958
rect 898 924 954 958
rect 988 924 1044 958
rect 1078 924 1137 958
rect 443 900 1137 924
rect 443 868 516 900
rect 550 868 616 900
rect 650 868 716 900
rect 750 868 816 900
rect 443 834 504 868
rect 550 866 594 868
rect 650 866 684 868
rect 750 866 774 868
rect 538 834 594 866
rect 628 834 684 866
rect 718 834 774 866
rect 808 866 816 868
rect 850 868 916 900
rect 850 866 864 868
rect 808 834 864 866
rect 898 866 916 868
rect 950 868 1016 900
rect 1050 868 1137 900
rect 950 866 954 868
rect 898 834 954 866
rect 988 866 1016 868
rect 988 834 1044 866
rect 1078 834 1137 868
rect 443 800 1137 834
rect 443 778 516 800
rect 550 778 616 800
rect 650 778 716 800
rect 750 778 816 800
rect 443 744 504 778
rect 550 766 594 778
rect 650 766 684 778
rect 750 766 774 778
rect 538 744 594 766
rect 628 744 684 766
rect 718 744 774 766
rect 808 766 816 778
rect 850 778 916 800
rect 850 766 864 778
rect 808 744 864 766
rect 898 766 916 778
rect 950 778 1016 800
rect 1050 778 1137 800
rect 950 766 954 778
rect 898 744 954 766
rect 988 766 1016 778
rect 988 744 1044 766
rect 1078 744 1137 778
rect 443 700 1137 744
rect 443 688 516 700
rect 550 688 616 700
rect 650 688 716 700
rect 750 688 816 700
rect 443 654 504 688
rect 550 666 594 688
rect 650 666 684 688
rect 750 666 774 688
rect 538 654 594 666
rect 628 654 684 666
rect 718 654 774 666
rect 808 666 816 688
rect 850 688 916 700
rect 850 666 864 688
rect 808 654 864 666
rect 898 666 916 688
rect 950 688 1016 700
rect 1050 688 1137 700
rect 950 666 954 688
rect 898 654 954 666
rect 988 666 1016 688
rect 988 654 1044 666
rect 1078 654 1137 688
rect 443 593 1137 654
rect 1199 1236 1271 1292
rect 1199 1202 1218 1236
rect 1252 1202 1271 1236
rect 1199 1146 1271 1202
rect 1199 1112 1218 1146
rect 1252 1112 1271 1146
rect 1199 1056 1271 1112
rect 1199 1022 1218 1056
rect 1252 1022 1271 1056
rect 1199 966 1271 1022
rect 1199 932 1218 966
rect 1252 932 1271 966
rect 1199 876 1271 932
rect 1199 842 1218 876
rect 1252 842 1271 876
rect 1199 786 1271 842
rect 1199 752 1218 786
rect 1252 752 1271 786
rect 1199 696 1271 752
rect 1199 662 1218 696
rect 1252 662 1271 696
rect 1199 606 1271 662
rect 309 531 381 591
rect 1199 572 1218 606
rect 1252 572 1271 606
rect 1199 531 1271 572
rect 309 512 1271 531
rect 309 478 406 512
rect 440 478 496 512
rect 530 478 586 512
rect 620 478 676 512
rect 710 478 766 512
rect 800 478 856 512
rect 890 478 946 512
rect 980 478 1036 512
rect 1070 478 1126 512
rect 1160 478 1271 512
rect 309 459 1271 478
rect 1335 1402 1367 1436
rect 1401 1402 1434 1436
rect 1335 1346 1434 1402
rect 1335 1312 1367 1346
rect 1401 1312 1434 1346
rect 1335 1256 1434 1312
rect 1335 1222 1367 1256
rect 1401 1222 1434 1256
rect 1335 1166 1434 1222
rect 1335 1132 1367 1166
rect 1401 1132 1434 1166
rect 1335 1076 1434 1132
rect 1335 1042 1367 1076
rect 1401 1042 1434 1076
rect 1335 986 1434 1042
rect 1335 952 1367 986
rect 1401 952 1434 986
rect 1335 896 1434 952
rect 1335 862 1367 896
rect 1401 862 1434 896
rect 1335 806 1434 862
rect 1335 772 1367 806
rect 1401 772 1434 806
rect 1335 716 1434 772
rect 1335 682 1367 716
rect 1401 682 1434 716
rect 1335 626 1434 682
rect 1335 592 1367 626
rect 1401 592 1434 626
rect 1335 536 1434 592
rect 1335 502 1367 536
rect 1401 502 1434 536
rect 146 412 180 446
rect 214 412 245 446
rect 146 395 245 412
rect 1335 446 1434 502
rect 1335 412 1367 446
rect 1401 412 1434 446
rect 1335 395 1434 412
rect 146 362 1434 395
rect 146 328 276 362
rect 310 328 366 362
rect 400 328 456 362
rect 490 328 546 362
rect 580 328 636 362
rect 670 328 726 362
rect 760 328 816 362
rect 850 328 906 362
rect 940 328 996 362
rect 1030 328 1086 362
rect 1120 328 1176 362
rect 1210 328 1266 362
rect 1300 328 1434 362
rect 146 296 1434 328
rect 120 17 1460 30
rect 120 -17 303 17
rect 337 -17 503 17
rect 537 -17 703 17
rect 737 -17 903 17
rect 937 -17 1103 17
rect 1137 -17 1303 17
rect 1337 -17 1460 17
rect 120 -30 1460 -17
<< viali >>
rect 303 1863 337 1897
rect 503 1863 537 1897
rect 703 1863 737 1897
rect 903 1863 937 1897
rect 1103 1863 1137 1897
rect 1303 1863 1337 1897
rect 516 1194 538 1200
rect 538 1194 550 1200
rect 616 1194 628 1200
rect 628 1194 650 1200
rect 716 1194 718 1200
rect 718 1194 750 1200
rect 516 1166 550 1194
rect 616 1166 650 1194
rect 716 1166 750 1194
rect 816 1166 850 1200
rect 916 1166 950 1200
rect 1016 1194 1044 1200
rect 1044 1194 1050 1200
rect 1016 1166 1050 1194
rect 516 1066 550 1100
rect 616 1066 650 1100
rect 716 1066 750 1100
rect 816 1066 850 1100
rect 916 1066 950 1100
rect 1016 1066 1050 1100
rect 516 966 550 1000
rect 616 966 650 1000
rect 716 966 750 1000
rect 816 966 850 1000
rect 916 966 950 1000
rect 1016 966 1050 1000
rect 516 868 550 900
rect 616 868 650 900
rect 716 868 750 900
rect 516 866 538 868
rect 538 866 550 868
rect 616 866 628 868
rect 628 866 650 868
rect 716 866 718 868
rect 718 866 750 868
rect 816 866 850 900
rect 916 866 950 900
rect 1016 868 1050 900
rect 1016 866 1044 868
rect 1044 866 1050 868
rect 516 778 550 800
rect 616 778 650 800
rect 716 778 750 800
rect 516 766 538 778
rect 538 766 550 778
rect 616 766 628 778
rect 628 766 650 778
rect 716 766 718 778
rect 718 766 750 778
rect 816 766 850 800
rect 916 766 950 800
rect 1016 778 1050 800
rect 1016 766 1044 778
rect 1044 766 1050 778
rect 516 688 550 700
rect 616 688 650 700
rect 716 688 750 700
rect 516 666 538 688
rect 538 666 550 688
rect 616 666 628 688
rect 628 666 650 688
rect 716 666 718 688
rect 718 666 750 688
rect 816 666 850 700
rect 916 666 950 700
rect 1016 688 1050 700
rect 1016 666 1044 688
rect 1044 666 1050 688
rect 303 -17 337 17
rect 503 -17 537 17
rect 703 -17 737 17
rect 903 -17 937 17
rect 1103 -17 1137 17
rect 1303 -17 1337 17
<< metal1 >>
rect 120 1897 1460 1940
rect 120 1863 303 1897
rect 337 1863 503 1897
rect 537 1863 703 1897
rect 737 1863 903 1897
rect 937 1863 1103 1897
rect 1137 1863 1303 1897
rect 1337 1863 1460 1897
rect 120 1820 1460 1863
rect 485 1200 1095 1245
rect 485 1166 516 1200
rect 550 1166 616 1200
rect 650 1166 716 1200
rect 750 1166 816 1200
rect 850 1166 916 1200
rect 950 1166 1016 1200
rect 1050 1166 1095 1200
rect 485 1100 1095 1166
rect 485 1066 516 1100
rect 550 1066 616 1100
rect 650 1066 716 1100
rect 750 1066 816 1100
rect 850 1066 916 1100
rect 950 1066 1016 1100
rect 1050 1066 1095 1100
rect 485 1000 1095 1066
rect 485 966 516 1000
rect 550 966 616 1000
rect 650 966 716 1000
rect 750 966 816 1000
rect 850 966 916 1000
rect 950 966 1016 1000
rect 1050 966 1095 1000
rect 485 900 1095 966
rect 485 866 516 900
rect 550 866 616 900
rect 650 866 716 900
rect 750 866 816 900
rect 850 866 916 900
rect 950 866 1016 900
rect 1050 866 1095 900
rect 485 800 1095 866
rect 485 766 516 800
rect 550 766 616 800
rect 650 766 716 800
rect 750 766 816 800
rect 850 766 916 800
rect 950 766 1016 800
rect 1050 766 1095 800
rect 485 700 1095 766
rect 485 666 516 700
rect 550 666 616 700
rect 650 666 716 700
rect 750 666 816 700
rect 850 666 916 700
rect 950 666 1016 700
rect 1050 666 1095 700
rect 485 635 1095 666
rect 120 17 1460 60
rect 120 -17 303 17
rect 337 -17 503 17
rect 537 -17 703 17
rect 737 -17 903 17
rect 937 -17 1103 17
rect 1137 -17 1303 17
rect 1337 -17 1460 17
rect 120 -60 1460 -17
<< labels >>
flabel locali s 674 896 922 1000 0 FreeSans 625 0 0 0 xm1/Emitter
port 1 nsew
flabel locali s 733 1522 834 1571 0 FreeSans 625 0 0 0 xm1/Collector
port 2 nsew
flabel locali s 710 1372 828 1412 0 FreeSans 625 0 0 0 xm1/Base
port 3 nsew
flabel locali s 682 1010 910 1140 1 FreeSans 750 0 0 0 Emitter
port 4 nsew
flabel locali s 894 1372 1014 1412 1 FreeSans 750 0 0 0 Base
port 5 nsew
flabel locali s 930 1524 1050 1564 1 FreeSans 750 0 0 0 Collector
port 6 nsew
flabel metal1 s 120 1850 180 1910 1 FreeSans 1250 0 0 0 VPWR
port 7 nsew
flabel metal1 s 120 -30 180 30 1 FreeSans 1250 0 0 0 VGND
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 1580 1880
<< end >>
