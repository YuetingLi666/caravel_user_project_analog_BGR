magic
tech sky130A
magscale 1 2
timestamp 1654901230
<< pwell >>
rect 120 1457 10840 1610
rect 120 423 273 1457
rect 1307 423 1613 1457
rect 2647 423 2953 1457
rect 3987 423 4293 1457
rect 5327 423 5633 1457
rect 6667 423 6973 1457
rect 8007 423 8313 1457
rect 9347 423 9653 1457
rect 10687 423 10840 1457
rect 120 270 10840 423
<< nbase >>
rect 273 423 1307 1457
rect 1613 423 2647 1457
rect 2953 423 3987 1457
rect 4293 423 5327 1457
rect 5633 423 6667 1457
rect 6973 423 8007 1457
rect 8313 423 9347 1457
rect 9653 423 10687 1457
<< pdiff >>
rect 450 1228 1130 1280
rect 450 1194 504 1228
rect 538 1194 594 1228
rect 628 1194 684 1228
rect 718 1194 774 1228
rect 808 1194 864 1228
rect 898 1194 954 1228
rect 988 1194 1044 1228
rect 1078 1194 1130 1228
rect 450 1138 1130 1194
rect 450 1104 504 1138
rect 538 1104 594 1138
rect 628 1104 684 1138
rect 718 1104 774 1138
rect 808 1104 864 1138
rect 898 1104 954 1138
rect 988 1104 1044 1138
rect 1078 1104 1130 1138
rect 450 1048 1130 1104
rect 450 1014 504 1048
rect 538 1014 594 1048
rect 628 1014 684 1048
rect 718 1014 774 1048
rect 808 1014 864 1048
rect 898 1014 954 1048
rect 988 1014 1044 1048
rect 1078 1014 1130 1048
rect 450 958 1130 1014
rect 450 924 504 958
rect 538 924 594 958
rect 628 924 684 958
rect 718 924 774 958
rect 808 924 864 958
rect 898 924 954 958
rect 988 924 1044 958
rect 1078 924 1130 958
rect 450 868 1130 924
rect 450 834 504 868
rect 538 834 594 868
rect 628 834 684 868
rect 718 834 774 868
rect 808 834 864 868
rect 898 834 954 868
rect 988 834 1044 868
rect 1078 834 1130 868
rect 450 778 1130 834
rect 450 744 504 778
rect 538 744 594 778
rect 628 744 684 778
rect 718 744 774 778
rect 808 744 864 778
rect 898 744 954 778
rect 988 744 1044 778
rect 1078 744 1130 778
rect 450 688 1130 744
rect 450 654 504 688
rect 538 654 594 688
rect 628 654 684 688
rect 718 654 774 688
rect 808 654 864 688
rect 898 654 954 688
rect 988 654 1044 688
rect 1078 654 1130 688
rect 450 600 1130 654
rect 1790 1228 2470 1280
rect 1790 1194 1844 1228
rect 1878 1194 1934 1228
rect 1968 1194 2024 1228
rect 2058 1194 2114 1228
rect 2148 1194 2204 1228
rect 2238 1194 2294 1228
rect 2328 1194 2384 1228
rect 2418 1194 2470 1228
rect 1790 1138 2470 1194
rect 1790 1104 1844 1138
rect 1878 1104 1934 1138
rect 1968 1104 2024 1138
rect 2058 1104 2114 1138
rect 2148 1104 2204 1138
rect 2238 1104 2294 1138
rect 2328 1104 2384 1138
rect 2418 1104 2470 1138
rect 1790 1048 2470 1104
rect 1790 1014 1844 1048
rect 1878 1014 1934 1048
rect 1968 1014 2024 1048
rect 2058 1014 2114 1048
rect 2148 1014 2204 1048
rect 2238 1014 2294 1048
rect 2328 1014 2384 1048
rect 2418 1014 2470 1048
rect 1790 958 2470 1014
rect 1790 924 1844 958
rect 1878 924 1934 958
rect 1968 924 2024 958
rect 2058 924 2114 958
rect 2148 924 2204 958
rect 2238 924 2294 958
rect 2328 924 2384 958
rect 2418 924 2470 958
rect 1790 868 2470 924
rect 1790 834 1844 868
rect 1878 834 1934 868
rect 1968 834 2024 868
rect 2058 834 2114 868
rect 2148 834 2204 868
rect 2238 834 2294 868
rect 2328 834 2384 868
rect 2418 834 2470 868
rect 1790 778 2470 834
rect 1790 744 1844 778
rect 1878 744 1934 778
rect 1968 744 2024 778
rect 2058 744 2114 778
rect 2148 744 2204 778
rect 2238 744 2294 778
rect 2328 744 2384 778
rect 2418 744 2470 778
rect 1790 688 2470 744
rect 1790 654 1844 688
rect 1878 654 1934 688
rect 1968 654 2024 688
rect 2058 654 2114 688
rect 2148 654 2204 688
rect 2238 654 2294 688
rect 2328 654 2384 688
rect 2418 654 2470 688
rect 1790 600 2470 654
rect 3130 1228 3810 1280
rect 3130 1194 3184 1228
rect 3218 1194 3274 1228
rect 3308 1194 3364 1228
rect 3398 1194 3454 1228
rect 3488 1194 3544 1228
rect 3578 1194 3634 1228
rect 3668 1194 3724 1228
rect 3758 1194 3810 1228
rect 3130 1138 3810 1194
rect 3130 1104 3184 1138
rect 3218 1104 3274 1138
rect 3308 1104 3364 1138
rect 3398 1104 3454 1138
rect 3488 1104 3544 1138
rect 3578 1104 3634 1138
rect 3668 1104 3724 1138
rect 3758 1104 3810 1138
rect 3130 1048 3810 1104
rect 3130 1014 3184 1048
rect 3218 1014 3274 1048
rect 3308 1014 3364 1048
rect 3398 1014 3454 1048
rect 3488 1014 3544 1048
rect 3578 1014 3634 1048
rect 3668 1014 3724 1048
rect 3758 1014 3810 1048
rect 3130 958 3810 1014
rect 3130 924 3184 958
rect 3218 924 3274 958
rect 3308 924 3364 958
rect 3398 924 3454 958
rect 3488 924 3544 958
rect 3578 924 3634 958
rect 3668 924 3724 958
rect 3758 924 3810 958
rect 3130 868 3810 924
rect 3130 834 3184 868
rect 3218 834 3274 868
rect 3308 834 3364 868
rect 3398 834 3454 868
rect 3488 834 3544 868
rect 3578 834 3634 868
rect 3668 834 3724 868
rect 3758 834 3810 868
rect 3130 778 3810 834
rect 3130 744 3184 778
rect 3218 744 3274 778
rect 3308 744 3364 778
rect 3398 744 3454 778
rect 3488 744 3544 778
rect 3578 744 3634 778
rect 3668 744 3724 778
rect 3758 744 3810 778
rect 3130 688 3810 744
rect 3130 654 3184 688
rect 3218 654 3274 688
rect 3308 654 3364 688
rect 3398 654 3454 688
rect 3488 654 3544 688
rect 3578 654 3634 688
rect 3668 654 3724 688
rect 3758 654 3810 688
rect 3130 600 3810 654
rect 4470 1228 5150 1280
rect 4470 1194 4524 1228
rect 4558 1194 4614 1228
rect 4648 1194 4704 1228
rect 4738 1194 4794 1228
rect 4828 1194 4884 1228
rect 4918 1194 4974 1228
rect 5008 1194 5064 1228
rect 5098 1194 5150 1228
rect 4470 1138 5150 1194
rect 4470 1104 4524 1138
rect 4558 1104 4614 1138
rect 4648 1104 4704 1138
rect 4738 1104 4794 1138
rect 4828 1104 4884 1138
rect 4918 1104 4974 1138
rect 5008 1104 5064 1138
rect 5098 1104 5150 1138
rect 4470 1048 5150 1104
rect 4470 1014 4524 1048
rect 4558 1014 4614 1048
rect 4648 1014 4704 1048
rect 4738 1014 4794 1048
rect 4828 1014 4884 1048
rect 4918 1014 4974 1048
rect 5008 1014 5064 1048
rect 5098 1014 5150 1048
rect 4470 958 5150 1014
rect 4470 924 4524 958
rect 4558 924 4614 958
rect 4648 924 4704 958
rect 4738 924 4794 958
rect 4828 924 4884 958
rect 4918 924 4974 958
rect 5008 924 5064 958
rect 5098 924 5150 958
rect 4470 868 5150 924
rect 4470 834 4524 868
rect 4558 834 4614 868
rect 4648 834 4704 868
rect 4738 834 4794 868
rect 4828 834 4884 868
rect 4918 834 4974 868
rect 5008 834 5064 868
rect 5098 834 5150 868
rect 4470 778 5150 834
rect 4470 744 4524 778
rect 4558 744 4614 778
rect 4648 744 4704 778
rect 4738 744 4794 778
rect 4828 744 4884 778
rect 4918 744 4974 778
rect 5008 744 5064 778
rect 5098 744 5150 778
rect 4470 688 5150 744
rect 4470 654 4524 688
rect 4558 654 4614 688
rect 4648 654 4704 688
rect 4738 654 4794 688
rect 4828 654 4884 688
rect 4918 654 4974 688
rect 5008 654 5064 688
rect 5098 654 5150 688
rect 4470 600 5150 654
rect 5810 1228 6490 1280
rect 5810 1194 5864 1228
rect 5898 1194 5954 1228
rect 5988 1194 6044 1228
rect 6078 1194 6134 1228
rect 6168 1194 6224 1228
rect 6258 1194 6314 1228
rect 6348 1194 6404 1228
rect 6438 1194 6490 1228
rect 5810 1138 6490 1194
rect 5810 1104 5864 1138
rect 5898 1104 5954 1138
rect 5988 1104 6044 1138
rect 6078 1104 6134 1138
rect 6168 1104 6224 1138
rect 6258 1104 6314 1138
rect 6348 1104 6404 1138
rect 6438 1104 6490 1138
rect 5810 1048 6490 1104
rect 5810 1014 5864 1048
rect 5898 1014 5954 1048
rect 5988 1014 6044 1048
rect 6078 1014 6134 1048
rect 6168 1014 6224 1048
rect 6258 1014 6314 1048
rect 6348 1014 6404 1048
rect 6438 1014 6490 1048
rect 5810 958 6490 1014
rect 5810 924 5864 958
rect 5898 924 5954 958
rect 5988 924 6044 958
rect 6078 924 6134 958
rect 6168 924 6224 958
rect 6258 924 6314 958
rect 6348 924 6404 958
rect 6438 924 6490 958
rect 5810 868 6490 924
rect 5810 834 5864 868
rect 5898 834 5954 868
rect 5988 834 6044 868
rect 6078 834 6134 868
rect 6168 834 6224 868
rect 6258 834 6314 868
rect 6348 834 6404 868
rect 6438 834 6490 868
rect 5810 778 6490 834
rect 5810 744 5864 778
rect 5898 744 5954 778
rect 5988 744 6044 778
rect 6078 744 6134 778
rect 6168 744 6224 778
rect 6258 744 6314 778
rect 6348 744 6404 778
rect 6438 744 6490 778
rect 5810 688 6490 744
rect 5810 654 5864 688
rect 5898 654 5954 688
rect 5988 654 6044 688
rect 6078 654 6134 688
rect 6168 654 6224 688
rect 6258 654 6314 688
rect 6348 654 6404 688
rect 6438 654 6490 688
rect 5810 600 6490 654
rect 7150 1228 7830 1280
rect 7150 1194 7204 1228
rect 7238 1194 7294 1228
rect 7328 1194 7384 1228
rect 7418 1194 7474 1228
rect 7508 1194 7564 1228
rect 7598 1194 7654 1228
rect 7688 1194 7744 1228
rect 7778 1194 7830 1228
rect 7150 1138 7830 1194
rect 7150 1104 7204 1138
rect 7238 1104 7294 1138
rect 7328 1104 7384 1138
rect 7418 1104 7474 1138
rect 7508 1104 7564 1138
rect 7598 1104 7654 1138
rect 7688 1104 7744 1138
rect 7778 1104 7830 1138
rect 7150 1048 7830 1104
rect 7150 1014 7204 1048
rect 7238 1014 7294 1048
rect 7328 1014 7384 1048
rect 7418 1014 7474 1048
rect 7508 1014 7564 1048
rect 7598 1014 7654 1048
rect 7688 1014 7744 1048
rect 7778 1014 7830 1048
rect 7150 958 7830 1014
rect 7150 924 7204 958
rect 7238 924 7294 958
rect 7328 924 7384 958
rect 7418 924 7474 958
rect 7508 924 7564 958
rect 7598 924 7654 958
rect 7688 924 7744 958
rect 7778 924 7830 958
rect 7150 868 7830 924
rect 7150 834 7204 868
rect 7238 834 7294 868
rect 7328 834 7384 868
rect 7418 834 7474 868
rect 7508 834 7564 868
rect 7598 834 7654 868
rect 7688 834 7744 868
rect 7778 834 7830 868
rect 7150 778 7830 834
rect 7150 744 7204 778
rect 7238 744 7294 778
rect 7328 744 7384 778
rect 7418 744 7474 778
rect 7508 744 7564 778
rect 7598 744 7654 778
rect 7688 744 7744 778
rect 7778 744 7830 778
rect 7150 688 7830 744
rect 7150 654 7204 688
rect 7238 654 7294 688
rect 7328 654 7384 688
rect 7418 654 7474 688
rect 7508 654 7564 688
rect 7598 654 7654 688
rect 7688 654 7744 688
rect 7778 654 7830 688
rect 7150 600 7830 654
rect 8490 1228 9170 1280
rect 8490 1194 8544 1228
rect 8578 1194 8634 1228
rect 8668 1194 8724 1228
rect 8758 1194 8814 1228
rect 8848 1194 8904 1228
rect 8938 1194 8994 1228
rect 9028 1194 9084 1228
rect 9118 1194 9170 1228
rect 8490 1138 9170 1194
rect 8490 1104 8544 1138
rect 8578 1104 8634 1138
rect 8668 1104 8724 1138
rect 8758 1104 8814 1138
rect 8848 1104 8904 1138
rect 8938 1104 8994 1138
rect 9028 1104 9084 1138
rect 9118 1104 9170 1138
rect 8490 1048 9170 1104
rect 8490 1014 8544 1048
rect 8578 1014 8634 1048
rect 8668 1014 8724 1048
rect 8758 1014 8814 1048
rect 8848 1014 8904 1048
rect 8938 1014 8994 1048
rect 9028 1014 9084 1048
rect 9118 1014 9170 1048
rect 8490 958 9170 1014
rect 8490 924 8544 958
rect 8578 924 8634 958
rect 8668 924 8724 958
rect 8758 924 8814 958
rect 8848 924 8904 958
rect 8938 924 8994 958
rect 9028 924 9084 958
rect 9118 924 9170 958
rect 8490 868 9170 924
rect 8490 834 8544 868
rect 8578 834 8634 868
rect 8668 834 8724 868
rect 8758 834 8814 868
rect 8848 834 8904 868
rect 8938 834 8994 868
rect 9028 834 9084 868
rect 9118 834 9170 868
rect 8490 778 9170 834
rect 8490 744 8544 778
rect 8578 744 8634 778
rect 8668 744 8724 778
rect 8758 744 8814 778
rect 8848 744 8904 778
rect 8938 744 8994 778
rect 9028 744 9084 778
rect 9118 744 9170 778
rect 8490 688 9170 744
rect 8490 654 8544 688
rect 8578 654 8634 688
rect 8668 654 8724 688
rect 8758 654 8814 688
rect 8848 654 8904 688
rect 8938 654 8994 688
rect 9028 654 9084 688
rect 9118 654 9170 688
rect 8490 600 9170 654
rect 9830 1228 10510 1280
rect 9830 1194 9884 1228
rect 9918 1194 9974 1228
rect 10008 1194 10064 1228
rect 10098 1194 10154 1228
rect 10188 1194 10244 1228
rect 10278 1194 10334 1228
rect 10368 1194 10424 1228
rect 10458 1194 10510 1228
rect 9830 1138 10510 1194
rect 9830 1104 9884 1138
rect 9918 1104 9974 1138
rect 10008 1104 10064 1138
rect 10098 1104 10154 1138
rect 10188 1104 10244 1138
rect 10278 1104 10334 1138
rect 10368 1104 10424 1138
rect 10458 1104 10510 1138
rect 9830 1048 10510 1104
rect 9830 1014 9884 1048
rect 9918 1014 9974 1048
rect 10008 1014 10064 1048
rect 10098 1014 10154 1048
rect 10188 1014 10244 1048
rect 10278 1014 10334 1048
rect 10368 1014 10424 1048
rect 10458 1014 10510 1048
rect 9830 958 10510 1014
rect 9830 924 9884 958
rect 9918 924 9974 958
rect 10008 924 10064 958
rect 10098 924 10154 958
rect 10188 924 10244 958
rect 10278 924 10334 958
rect 10368 924 10424 958
rect 10458 924 10510 958
rect 9830 868 10510 924
rect 9830 834 9884 868
rect 9918 834 9974 868
rect 10008 834 10064 868
rect 10098 834 10154 868
rect 10188 834 10244 868
rect 10278 834 10334 868
rect 10368 834 10424 868
rect 10458 834 10510 868
rect 9830 778 10510 834
rect 9830 744 9884 778
rect 9918 744 9974 778
rect 10008 744 10064 778
rect 10098 744 10154 778
rect 10188 744 10244 778
rect 10278 744 10334 778
rect 10368 744 10424 778
rect 10458 744 10510 778
rect 9830 688 10510 744
rect 9830 654 9884 688
rect 9918 654 9974 688
rect 10008 654 10064 688
rect 10098 654 10154 688
rect 10188 654 10244 688
rect 10278 654 10334 688
rect 10368 654 10424 688
rect 10458 654 10510 688
rect 9830 600 10510 654
<< pdiffc >>
rect 504 1194 538 1228
rect 594 1194 628 1228
rect 684 1194 718 1228
rect 774 1194 808 1228
rect 864 1194 898 1228
rect 954 1194 988 1228
rect 1044 1194 1078 1228
rect 504 1104 538 1138
rect 594 1104 628 1138
rect 684 1104 718 1138
rect 774 1104 808 1138
rect 864 1104 898 1138
rect 954 1104 988 1138
rect 1044 1104 1078 1138
rect 504 1014 538 1048
rect 594 1014 628 1048
rect 684 1014 718 1048
rect 774 1014 808 1048
rect 864 1014 898 1048
rect 954 1014 988 1048
rect 1044 1014 1078 1048
rect 504 924 538 958
rect 594 924 628 958
rect 684 924 718 958
rect 774 924 808 958
rect 864 924 898 958
rect 954 924 988 958
rect 1044 924 1078 958
rect 504 834 538 868
rect 594 834 628 868
rect 684 834 718 868
rect 774 834 808 868
rect 864 834 898 868
rect 954 834 988 868
rect 1044 834 1078 868
rect 504 744 538 778
rect 594 744 628 778
rect 684 744 718 778
rect 774 744 808 778
rect 864 744 898 778
rect 954 744 988 778
rect 1044 744 1078 778
rect 504 654 538 688
rect 594 654 628 688
rect 684 654 718 688
rect 774 654 808 688
rect 864 654 898 688
rect 954 654 988 688
rect 1044 654 1078 688
rect 1844 1194 1878 1228
rect 1934 1194 1968 1228
rect 2024 1194 2058 1228
rect 2114 1194 2148 1228
rect 2204 1194 2238 1228
rect 2294 1194 2328 1228
rect 2384 1194 2418 1228
rect 1844 1104 1878 1138
rect 1934 1104 1968 1138
rect 2024 1104 2058 1138
rect 2114 1104 2148 1138
rect 2204 1104 2238 1138
rect 2294 1104 2328 1138
rect 2384 1104 2418 1138
rect 1844 1014 1878 1048
rect 1934 1014 1968 1048
rect 2024 1014 2058 1048
rect 2114 1014 2148 1048
rect 2204 1014 2238 1048
rect 2294 1014 2328 1048
rect 2384 1014 2418 1048
rect 1844 924 1878 958
rect 1934 924 1968 958
rect 2024 924 2058 958
rect 2114 924 2148 958
rect 2204 924 2238 958
rect 2294 924 2328 958
rect 2384 924 2418 958
rect 1844 834 1878 868
rect 1934 834 1968 868
rect 2024 834 2058 868
rect 2114 834 2148 868
rect 2204 834 2238 868
rect 2294 834 2328 868
rect 2384 834 2418 868
rect 1844 744 1878 778
rect 1934 744 1968 778
rect 2024 744 2058 778
rect 2114 744 2148 778
rect 2204 744 2238 778
rect 2294 744 2328 778
rect 2384 744 2418 778
rect 1844 654 1878 688
rect 1934 654 1968 688
rect 2024 654 2058 688
rect 2114 654 2148 688
rect 2204 654 2238 688
rect 2294 654 2328 688
rect 2384 654 2418 688
rect 3184 1194 3218 1228
rect 3274 1194 3308 1228
rect 3364 1194 3398 1228
rect 3454 1194 3488 1228
rect 3544 1194 3578 1228
rect 3634 1194 3668 1228
rect 3724 1194 3758 1228
rect 3184 1104 3218 1138
rect 3274 1104 3308 1138
rect 3364 1104 3398 1138
rect 3454 1104 3488 1138
rect 3544 1104 3578 1138
rect 3634 1104 3668 1138
rect 3724 1104 3758 1138
rect 3184 1014 3218 1048
rect 3274 1014 3308 1048
rect 3364 1014 3398 1048
rect 3454 1014 3488 1048
rect 3544 1014 3578 1048
rect 3634 1014 3668 1048
rect 3724 1014 3758 1048
rect 3184 924 3218 958
rect 3274 924 3308 958
rect 3364 924 3398 958
rect 3454 924 3488 958
rect 3544 924 3578 958
rect 3634 924 3668 958
rect 3724 924 3758 958
rect 3184 834 3218 868
rect 3274 834 3308 868
rect 3364 834 3398 868
rect 3454 834 3488 868
rect 3544 834 3578 868
rect 3634 834 3668 868
rect 3724 834 3758 868
rect 3184 744 3218 778
rect 3274 744 3308 778
rect 3364 744 3398 778
rect 3454 744 3488 778
rect 3544 744 3578 778
rect 3634 744 3668 778
rect 3724 744 3758 778
rect 3184 654 3218 688
rect 3274 654 3308 688
rect 3364 654 3398 688
rect 3454 654 3488 688
rect 3544 654 3578 688
rect 3634 654 3668 688
rect 3724 654 3758 688
rect 4524 1194 4558 1228
rect 4614 1194 4648 1228
rect 4704 1194 4738 1228
rect 4794 1194 4828 1228
rect 4884 1194 4918 1228
rect 4974 1194 5008 1228
rect 5064 1194 5098 1228
rect 4524 1104 4558 1138
rect 4614 1104 4648 1138
rect 4704 1104 4738 1138
rect 4794 1104 4828 1138
rect 4884 1104 4918 1138
rect 4974 1104 5008 1138
rect 5064 1104 5098 1138
rect 4524 1014 4558 1048
rect 4614 1014 4648 1048
rect 4704 1014 4738 1048
rect 4794 1014 4828 1048
rect 4884 1014 4918 1048
rect 4974 1014 5008 1048
rect 5064 1014 5098 1048
rect 4524 924 4558 958
rect 4614 924 4648 958
rect 4704 924 4738 958
rect 4794 924 4828 958
rect 4884 924 4918 958
rect 4974 924 5008 958
rect 5064 924 5098 958
rect 4524 834 4558 868
rect 4614 834 4648 868
rect 4704 834 4738 868
rect 4794 834 4828 868
rect 4884 834 4918 868
rect 4974 834 5008 868
rect 5064 834 5098 868
rect 4524 744 4558 778
rect 4614 744 4648 778
rect 4704 744 4738 778
rect 4794 744 4828 778
rect 4884 744 4918 778
rect 4974 744 5008 778
rect 5064 744 5098 778
rect 4524 654 4558 688
rect 4614 654 4648 688
rect 4704 654 4738 688
rect 4794 654 4828 688
rect 4884 654 4918 688
rect 4974 654 5008 688
rect 5064 654 5098 688
rect 5864 1194 5898 1228
rect 5954 1194 5988 1228
rect 6044 1194 6078 1228
rect 6134 1194 6168 1228
rect 6224 1194 6258 1228
rect 6314 1194 6348 1228
rect 6404 1194 6438 1228
rect 5864 1104 5898 1138
rect 5954 1104 5988 1138
rect 6044 1104 6078 1138
rect 6134 1104 6168 1138
rect 6224 1104 6258 1138
rect 6314 1104 6348 1138
rect 6404 1104 6438 1138
rect 5864 1014 5898 1048
rect 5954 1014 5988 1048
rect 6044 1014 6078 1048
rect 6134 1014 6168 1048
rect 6224 1014 6258 1048
rect 6314 1014 6348 1048
rect 6404 1014 6438 1048
rect 5864 924 5898 958
rect 5954 924 5988 958
rect 6044 924 6078 958
rect 6134 924 6168 958
rect 6224 924 6258 958
rect 6314 924 6348 958
rect 6404 924 6438 958
rect 5864 834 5898 868
rect 5954 834 5988 868
rect 6044 834 6078 868
rect 6134 834 6168 868
rect 6224 834 6258 868
rect 6314 834 6348 868
rect 6404 834 6438 868
rect 5864 744 5898 778
rect 5954 744 5988 778
rect 6044 744 6078 778
rect 6134 744 6168 778
rect 6224 744 6258 778
rect 6314 744 6348 778
rect 6404 744 6438 778
rect 5864 654 5898 688
rect 5954 654 5988 688
rect 6044 654 6078 688
rect 6134 654 6168 688
rect 6224 654 6258 688
rect 6314 654 6348 688
rect 6404 654 6438 688
rect 7204 1194 7238 1228
rect 7294 1194 7328 1228
rect 7384 1194 7418 1228
rect 7474 1194 7508 1228
rect 7564 1194 7598 1228
rect 7654 1194 7688 1228
rect 7744 1194 7778 1228
rect 7204 1104 7238 1138
rect 7294 1104 7328 1138
rect 7384 1104 7418 1138
rect 7474 1104 7508 1138
rect 7564 1104 7598 1138
rect 7654 1104 7688 1138
rect 7744 1104 7778 1138
rect 7204 1014 7238 1048
rect 7294 1014 7328 1048
rect 7384 1014 7418 1048
rect 7474 1014 7508 1048
rect 7564 1014 7598 1048
rect 7654 1014 7688 1048
rect 7744 1014 7778 1048
rect 7204 924 7238 958
rect 7294 924 7328 958
rect 7384 924 7418 958
rect 7474 924 7508 958
rect 7564 924 7598 958
rect 7654 924 7688 958
rect 7744 924 7778 958
rect 7204 834 7238 868
rect 7294 834 7328 868
rect 7384 834 7418 868
rect 7474 834 7508 868
rect 7564 834 7598 868
rect 7654 834 7688 868
rect 7744 834 7778 868
rect 7204 744 7238 778
rect 7294 744 7328 778
rect 7384 744 7418 778
rect 7474 744 7508 778
rect 7564 744 7598 778
rect 7654 744 7688 778
rect 7744 744 7778 778
rect 7204 654 7238 688
rect 7294 654 7328 688
rect 7384 654 7418 688
rect 7474 654 7508 688
rect 7564 654 7598 688
rect 7654 654 7688 688
rect 7744 654 7778 688
rect 8544 1194 8578 1228
rect 8634 1194 8668 1228
rect 8724 1194 8758 1228
rect 8814 1194 8848 1228
rect 8904 1194 8938 1228
rect 8994 1194 9028 1228
rect 9084 1194 9118 1228
rect 8544 1104 8578 1138
rect 8634 1104 8668 1138
rect 8724 1104 8758 1138
rect 8814 1104 8848 1138
rect 8904 1104 8938 1138
rect 8994 1104 9028 1138
rect 9084 1104 9118 1138
rect 8544 1014 8578 1048
rect 8634 1014 8668 1048
rect 8724 1014 8758 1048
rect 8814 1014 8848 1048
rect 8904 1014 8938 1048
rect 8994 1014 9028 1048
rect 9084 1014 9118 1048
rect 8544 924 8578 958
rect 8634 924 8668 958
rect 8724 924 8758 958
rect 8814 924 8848 958
rect 8904 924 8938 958
rect 8994 924 9028 958
rect 9084 924 9118 958
rect 8544 834 8578 868
rect 8634 834 8668 868
rect 8724 834 8758 868
rect 8814 834 8848 868
rect 8904 834 8938 868
rect 8994 834 9028 868
rect 9084 834 9118 868
rect 8544 744 8578 778
rect 8634 744 8668 778
rect 8724 744 8758 778
rect 8814 744 8848 778
rect 8904 744 8938 778
rect 8994 744 9028 778
rect 9084 744 9118 778
rect 8544 654 8578 688
rect 8634 654 8668 688
rect 8724 654 8758 688
rect 8814 654 8848 688
rect 8904 654 8938 688
rect 8994 654 9028 688
rect 9084 654 9118 688
rect 9884 1194 9918 1228
rect 9974 1194 10008 1228
rect 10064 1194 10098 1228
rect 10154 1194 10188 1228
rect 10244 1194 10278 1228
rect 10334 1194 10368 1228
rect 10424 1194 10458 1228
rect 9884 1104 9918 1138
rect 9974 1104 10008 1138
rect 10064 1104 10098 1138
rect 10154 1104 10188 1138
rect 10244 1104 10278 1138
rect 10334 1104 10368 1138
rect 10424 1104 10458 1138
rect 9884 1014 9918 1048
rect 9974 1014 10008 1048
rect 10064 1014 10098 1048
rect 10154 1014 10188 1048
rect 10244 1014 10278 1048
rect 10334 1014 10368 1048
rect 10424 1014 10458 1048
rect 9884 924 9918 958
rect 9974 924 10008 958
rect 10064 924 10098 958
rect 10154 924 10188 958
rect 10244 924 10278 958
rect 10334 924 10368 958
rect 10424 924 10458 958
rect 9884 834 9918 868
rect 9974 834 10008 868
rect 10064 834 10098 868
rect 10154 834 10188 868
rect 10244 834 10278 868
rect 10334 834 10368 868
rect 10424 834 10458 868
rect 9884 744 9918 778
rect 9974 744 10008 778
rect 10064 744 10098 778
rect 10154 744 10188 778
rect 10244 744 10278 778
rect 10334 744 10368 778
rect 10424 744 10458 778
rect 9884 654 9918 688
rect 9974 654 10008 688
rect 10064 654 10098 688
rect 10154 654 10188 688
rect 10244 654 10278 688
rect 10334 654 10368 688
rect 10424 654 10458 688
<< psubdiff >>
rect 146 1549 10814 1584
rect 146 1526 276 1549
rect 146 1492 180 1526
rect 214 1515 276 1526
rect 310 1515 366 1549
rect 400 1515 456 1549
rect 490 1515 546 1549
rect 580 1515 636 1549
rect 670 1515 726 1549
rect 760 1515 816 1549
rect 850 1515 906 1549
rect 940 1515 996 1549
rect 1030 1515 1086 1549
rect 1120 1515 1176 1549
rect 1210 1515 1266 1549
rect 1300 1526 1616 1549
rect 1300 1515 1367 1526
rect 214 1492 1367 1515
rect 1401 1492 1520 1526
rect 1554 1515 1616 1526
rect 1650 1515 1706 1549
rect 1740 1515 1796 1549
rect 1830 1515 1886 1549
rect 1920 1515 1976 1549
rect 2010 1515 2066 1549
rect 2100 1515 2156 1549
rect 2190 1515 2246 1549
rect 2280 1515 2336 1549
rect 2370 1515 2426 1549
rect 2460 1515 2516 1549
rect 2550 1515 2606 1549
rect 2640 1526 2956 1549
rect 2640 1515 2707 1526
rect 1554 1492 2707 1515
rect 2741 1492 2860 1526
rect 2894 1515 2956 1526
rect 2990 1515 3046 1549
rect 3080 1515 3136 1549
rect 3170 1515 3226 1549
rect 3260 1515 3316 1549
rect 3350 1515 3406 1549
rect 3440 1515 3496 1549
rect 3530 1515 3586 1549
rect 3620 1515 3676 1549
rect 3710 1515 3766 1549
rect 3800 1515 3856 1549
rect 3890 1515 3946 1549
rect 3980 1526 4296 1549
rect 3980 1515 4047 1526
rect 2894 1492 4047 1515
rect 4081 1492 4200 1526
rect 4234 1515 4296 1526
rect 4330 1515 4386 1549
rect 4420 1515 4476 1549
rect 4510 1515 4566 1549
rect 4600 1515 4656 1549
rect 4690 1515 4746 1549
rect 4780 1515 4836 1549
rect 4870 1515 4926 1549
rect 4960 1515 5016 1549
rect 5050 1515 5106 1549
rect 5140 1515 5196 1549
rect 5230 1515 5286 1549
rect 5320 1526 5636 1549
rect 5320 1515 5387 1526
rect 4234 1492 5387 1515
rect 5421 1492 5540 1526
rect 5574 1515 5636 1526
rect 5670 1515 5726 1549
rect 5760 1515 5816 1549
rect 5850 1515 5906 1549
rect 5940 1515 5996 1549
rect 6030 1515 6086 1549
rect 6120 1515 6176 1549
rect 6210 1515 6266 1549
rect 6300 1515 6356 1549
rect 6390 1515 6446 1549
rect 6480 1515 6536 1549
rect 6570 1515 6626 1549
rect 6660 1526 6976 1549
rect 6660 1515 6727 1526
rect 5574 1492 6727 1515
rect 6761 1492 6880 1526
rect 6914 1515 6976 1526
rect 7010 1515 7066 1549
rect 7100 1515 7156 1549
rect 7190 1515 7246 1549
rect 7280 1515 7336 1549
rect 7370 1515 7426 1549
rect 7460 1515 7516 1549
rect 7550 1515 7606 1549
rect 7640 1515 7696 1549
rect 7730 1515 7786 1549
rect 7820 1515 7876 1549
rect 7910 1515 7966 1549
rect 8000 1526 8316 1549
rect 8000 1515 8067 1526
rect 6914 1492 8067 1515
rect 8101 1492 8220 1526
rect 8254 1515 8316 1526
rect 8350 1515 8406 1549
rect 8440 1515 8496 1549
rect 8530 1515 8586 1549
rect 8620 1515 8676 1549
rect 8710 1515 8766 1549
rect 8800 1515 8856 1549
rect 8890 1515 8946 1549
rect 8980 1515 9036 1549
rect 9070 1515 9126 1549
rect 9160 1515 9216 1549
rect 9250 1515 9306 1549
rect 9340 1526 9656 1549
rect 9340 1515 9407 1526
rect 8254 1492 9407 1515
rect 9441 1492 9560 1526
rect 9594 1515 9656 1526
rect 9690 1515 9746 1549
rect 9780 1515 9836 1549
rect 9870 1515 9926 1549
rect 9960 1515 10016 1549
rect 10050 1515 10106 1549
rect 10140 1515 10196 1549
rect 10230 1515 10286 1549
rect 10320 1515 10376 1549
rect 10410 1515 10466 1549
rect 10500 1515 10556 1549
rect 10590 1515 10646 1549
rect 10680 1526 10814 1549
rect 10680 1515 10747 1526
rect 9594 1492 10747 1515
rect 10781 1492 10814 1526
rect 146 1483 10814 1492
rect 146 1436 247 1483
rect 146 1402 180 1436
rect 214 1402 247 1436
rect 1333 1436 1587 1483
rect 146 1346 247 1402
rect 146 1312 180 1346
rect 214 1312 247 1346
rect 146 1256 247 1312
rect 146 1222 180 1256
rect 214 1222 247 1256
rect 146 1166 247 1222
rect 146 1132 180 1166
rect 214 1132 247 1166
rect 146 1076 247 1132
rect 146 1042 180 1076
rect 214 1042 247 1076
rect 146 986 247 1042
rect 146 952 180 986
rect 214 952 247 986
rect 146 896 247 952
rect 146 862 180 896
rect 214 862 247 896
rect 146 806 247 862
rect 146 772 180 806
rect 214 772 247 806
rect 146 716 247 772
rect 146 682 180 716
rect 214 682 247 716
rect 146 626 247 682
rect 146 592 180 626
rect 214 592 247 626
rect 146 536 247 592
rect 146 502 180 536
rect 214 502 247 536
rect 146 446 247 502
rect 1333 1402 1367 1436
rect 1401 1402 1520 1436
rect 1554 1402 1587 1436
rect 2673 1436 2927 1483
rect 1333 1346 1587 1402
rect 1333 1312 1367 1346
rect 1401 1312 1520 1346
rect 1554 1312 1587 1346
rect 1333 1256 1587 1312
rect 1333 1222 1367 1256
rect 1401 1222 1520 1256
rect 1554 1222 1587 1256
rect 1333 1166 1587 1222
rect 1333 1132 1367 1166
rect 1401 1132 1520 1166
rect 1554 1132 1587 1166
rect 1333 1076 1587 1132
rect 1333 1042 1367 1076
rect 1401 1042 1520 1076
rect 1554 1042 1587 1076
rect 1333 986 1587 1042
rect 1333 952 1367 986
rect 1401 952 1520 986
rect 1554 952 1587 986
rect 1333 896 1587 952
rect 1333 862 1367 896
rect 1401 862 1520 896
rect 1554 862 1587 896
rect 1333 806 1587 862
rect 1333 772 1367 806
rect 1401 772 1520 806
rect 1554 772 1587 806
rect 1333 716 1587 772
rect 1333 682 1367 716
rect 1401 682 1520 716
rect 1554 682 1587 716
rect 1333 626 1587 682
rect 1333 592 1367 626
rect 1401 592 1520 626
rect 1554 592 1587 626
rect 1333 536 1587 592
rect 1333 502 1367 536
rect 1401 502 1520 536
rect 1554 502 1587 536
rect 146 412 180 446
rect 214 412 247 446
rect 146 397 247 412
rect 1333 446 1587 502
rect 2673 1402 2707 1436
rect 2741 1402 2860 1436
rect 2894 1402 2927 1436
rect 4013 1436 4267 1483
rect 2673 1346 2927 1402
rect 2673 1312 2707 1346
rect 2741 1312 2860 1346
rect 2894 1312 2927 1346
rect 2673 1256 2927 1312
rect 2673 1222 2707 1256
rect 2741 1222 2860 1256
rect 2894 1222 2927 1256
rect 2673 1166 2927 1222
rect 2673 1132 2707 1166
rect 2741 1132 2860 1166
rect 2894 1132 2927 1166
rect 2673 1076 2927 1132
rect 2673 1042 2707 1076
rect 2741 1042 2860 1076
rect 2894 1042 2927 1076
rect 2673 986 2927 1042
rect 2673 952 2707 986
rect 2741 952 2860 986
rect 2894 952 2927 986
rect 2673 896 2927 952
rect 2673 862 2707 896
rect 2741 862 2860 896
rect 2894 862 2927 896
rect 2673 806 2927 862
rect 2673 772 2707 806
rect 2741 772 2860 806
rect 2894 772 2927 806
rect 2673 716 2927 772
rect 2673 682 2707 716
rect 2741 682 2860 716
rect 2894 682 2927 716
rect 2673 626 2927 682
rect 2673 592 2707 626
rect 2741 592 2860 626
rect 2894 592 2927 626
rect 2673 536 2927 592
rect 2673 502 2707 536
rect 2741 502 2860 536
rect 2894 502 2927 536
rect 1333 412 1367 446
rect 1401 412 1520 446
rect 1554 412 1587 446
rect 1333 397 1587 412
rect 2673 446 2927 502
rect 4013 1402 4047 1436
rect 4081 1402 4200 1436
rect 4234 1402 4267 1436
rect 5353 1436 5607 1483
rect 4013 1346 4267 1402
rect 4013 1312 4047 1346
rect 4081 1312 4200 1346
rect 4234 1312 4267 1346
rect 4013 1256 4267 1312
rect 4013 1222 4047 1256
rect 4081 1222 4200 1256
rect 4234 1222 4267 1256
rect 4013 1166 4267 1222
rect 4013 1132 4047 1166
rect 4081 1132 4200 1166
rect 4234 1132 4267 1166
rect 4013 1076 4267 1132
rect 4013 1042 4047 1076
rect 4081 1042 4200 1076
rect 4234 1042 4267 1076
rect 4013 986 4267 1042
rect 4013 952 4047 986
rect 4081 952 4200 986
rect 4234 952 4267 986
rect 4013 896 4267 952
rect 4013 862 4047 896
rect 4081 862 4200 896
rect 4234 862 4267 896
rect 4013 806 4267 862
rect 4013 772 4047 806
rect 4081 772 4200 806
rect 4234 772 4267 806
rect 4013 716 4267 772
rect 4013 682 4047 716
rect 4081 682 4200 716
rect 4234 682 4267 716
rect 4013 626 4267 682
rect 4013 592 4047 626
rect 4081 592 4200 626
rect 4234 592 4267 626
rect 4013 536 4267 592
rect 4013 502 4047 536
rect 4081 502 4200 536
rect 4234 502 4267 536
rect 2673 412 2707 446
rect 2741 412 2860 446
rect 2894 412 2927 446
rect 2673 397 2927 412
rect 4013 446 4267 502
rect 5353 1402 5387 1436
rect 5421 1402 5540 1436
rect 5574 1402 5607 1436
rect 6693 1436 6947 1483
rect 5353 1346 5607 1402
rect 5353 1312 5387 1346
rect 5421 1312 5540 1346
rect 5574 1312 5607 1346
rect 5353 1256 5607 1312
rect 5353 1222 5387 1256
rect 5421 1222 5540 1256
rect 5574 1222 5607 1256
rect 5353 1166 5607 1222
rect 5353 1132 5387 1166
rect 5421 1132 5540 1166
rect 5574 1132 5607 1166
rect 5353 1076 5607 1132
rect 5353 1042 5387 1076
rect 5421 1042 5540 1076
rect 5574 1042 5607 1076
rect 5353 986 5607 1042
rect 5353 952 5387 986
rect 5421 952 5540 986
rect 5574 952 5607 986
rect 5353 896 5607 952
rect 5353 862 5387 896
rect 5421 862 5540 896
rect 5574 862 5607 896
rect 5353 806 5607 862
rect 5353 772 5387 806
rect 5421 772 5540 806
rect 5574 772 5607 806
rect 5353 716 5607 772
rect 5353 682 5387 716
rect 5421 682 5540 716
rect 5574 682 5607 716
rect 5353 626 5607 682
rect 5353 592 5387 626
rect 5421 592 5540 626
rect 5574 592 5607 626
rect 5353 536 5607 592
rect 5353 502 5387 536
rect 5421 502 5540 536
rect 5574 502 5607 536
rect 4013 412 4047 446
rect 4081 412 4200 446
rect 4234 412 4267 446
rect 4013 397 4267 412
rect 5353 446 5607 502
rect 6693 1402 6727 1436
rect 6761 1402 6880 1436
rect 6914 1402 6947 1436
rect 8033 1436 8287 1483
rect 6693 1346 6947 1402
rect 6693 1312 6727 1346
rect 6761 1312 6880 1346
rect 6914 1312 6947 1346
rect 6693 1256 6947 1312
rect 6693 1222 6727 1256
rect 6761 1222 6880 1256
rect 6914 1222 6947 1256
rect 6693 1166 6947 1222
rect 6693 1132 6727 1166
rect 6761 1132 6880 1166
rect 6914 1132 6947 1166
rect 6693 1076 6947 1132
rect 6693 1042 6727 1076
rect 6761 1042 6880 1076
rect 6914 1042 6947 1076
rect 6693 986 6947 1042
rect 6693 952 6727 986
rect 6761 952 6880 986
rect 6914 952 6947 986
rect 6693 896 6947 952
rect 6693 862 6727 896
rect 6761 862 6880 896
rect 6914 862 6947 896
rect 6693 806 6947 862
rect 6693 772 6727 806
rect 6761 772 6880 806
rect 6914 772 6947 806
rect 6693 716 6947 772
rect 6693 682 6727 716
rect 6761 682 6880 716
rect 6914 682 6947 716
rect 6693 626 6947 682
rect 6693 592 6727 626
rect 6761 592 6880 626
rect 6914 592 6947 626
rect 6693 536 6947 592
rect 6693 502 6727 536
rect 6761 502 6880 536
rect 6914 502 6947 536
rect 5353 412 5387 446
rect 5421 412 5540 446
rect 5574 412 5607 446
rect 5353 397 5607 412
rect 6693 446 6947 502
rect 8033 1402 8067 1436
rect 8101 1402 8220 1436
rect 8254 1402 8287 1436
rect 9373 1436 9627 1483
rect 8033 1346 8287 1402
rect 8033 1312 8067 1346
rect 8101 1312 8220 1346
rect 8254 1312 8287 1346
rect 8033 1256 8287 1312
rect 8033 1222 8067 1256
rect 8101 1222 8220 1256
rect 8254 1222 8287 1256
rect 8033 1166 8287 1222
rect 8033 1132 8067 1166
rect 8101 1132 8220 1166
rect 8254 1132 8287 1166
rect 8033 1076 8287 1132
rect 8033 1042 8067 1076
rect 8101 1042 8220 1076
rect 8254 1042 8287 1076
rect 8033 986 8287 1042
rect 8033 952 8067 986
rect 8101 952 8220 986
rect 8254 952 8287 986
rect 8033 896 8287 952
rect 8033 862 8067 896
rect 8101 862 8220 896
rect 8254 862 8287 896
rect 8033 806 8287 862
rect 8033 772 8067 806
rect 8101 772 8220 806
rect 8254 772 8287 806
rect 8033 716 8287 772
rect 8033 682 8067 716
rect 8101 682 8220 716
rect 8254 682 8287 716
rect 8033 626 8287 682
rect 8033 592 8067 626
rect 8101 592 8220 626
rect 8254 592 8287 626
rect 8033 536 8287 592
rect 8033 502 8067 536
rect 8101 502 8220 536
rect 8254 502 8287 536
rect 6693 412 6727 446
rect 6761 412 6880 446
rect 6914 412 6947 446
rect 6693 397 6947 412
rect 8033 446 8287 502
rect 9373 1402 9407 1436
rect 9441 1402 9560 1436
rect 9594 1402 9627 1436
rect 10713 1436 10814 1483
rect 9373 1346 9627 1402
rect 9373 1312 9407 1346
rect 9441 1312 9560 1346
rect 9594 1312 9627 1346
rect 9373 1256 9627 1312
rect 9373 1222 9407 1256
rect 9441 1222 9560 1256
rect 9594 1222 9627 1256
rect 9373 1166 9627 1222
rect 9373 1132 9407 1166
rect 9441 1132 9560 1166
rect 9594 1132 9627 1166
rect 9373 1076 9627 1132
rect 9373 1042 9407 1076
rect 9441 1042 9560 1076
rect 9594 1042 9627 1076
rect 9373 986 9627 1042
rect 9373 952 9407 986
rect 9441 952 9560 986
rect 9594 952 9627 986
rect 9373 896 9627 952
rect 9373 862 9407 896
rect 9441 862 9560 896
rect 9594 862 9627 896
rect 9373 806 9627 862
rect 9373 772 9407 806
rect 9441 772 9560 806
rect 9594 772 9627 806
rect 9373 716 9627 772
rect 9373 682 9407 716
rect 9441 682 9560 716
rect 9594 682 9627 716
rect 9373 626 9627 682
rect 9373 592 9407 626
rect 9441 592 9560 626
rect 9594 592 9627 626
rect 9373 536 9627 592
rect 9373 502 9407 536
rect 9441 502 9560 536
rect 9594 502 9627 536
rect 8033 412 8067 446
rect 8101 412 8220 446
rect 8254 412 8287 446
rect 8033 397 8287 412
rect 9373 446 9627 502
rect 10713 1402 10747 1436
rect 10781 1402 10814 1436
rect 10713 1346 10814 1402
rect 10713 1312 10747 1346
rect 10781 1312 10814 1346
rect 10713 1256 10814 1312
rect 10713 1222 10747 1256
rect 10781 1222 10814 1256
rect 10713 1166 10814 1222
rect 10713 1132 10747 1166
rect 10781 1132 10814 1166
rect 10713 1076 10814 1132
rect 10713 1042 10747 1076
rect 10781 1042 10814 1076
rect 10713 986 10814 1042
rect 10713 952 10747 986
rect 10781 952 10814 986
rect 10713 896 10814 952
rect 10713 862 10747 896
rect 10781 862 10814 896
rect 10713 806 10814 862
rect 10713 772 10747 806
rect 10781 772 10814 806
rect 10713 716 10814 772
rect 10713 682 10747 716
rect 10781 682 10814 716
rect 10713 626 10814 682
rect 10713 592 10747 626
rect 10781 592 10814 626
rect 10713 536 10814 592
rect 10713 502 10747 536
rect 10781 502 10814 536
rect 9373 412 9407 446
rect 9441 412 9560 446
rect 9594 412 9627 446
rect 9373 397 9627 412
rect 10713 446 10814 502
rect 10713 412 10747 446
rect 10781 412 10814 446
rect 10713 397 10814 412
rect 146 362 10814 397
rect 146 328 276 362
rect 310 328 366 362
rect 400 328 456 362
rect 490 328 546 362
rect 580 328 636 362
rect 670 328 726 362
rect 760 328 816 362
rect 850 328 906 362
rect 940 328 996 362
rect 1030 328 1086 362
rect 1120 328 1176 362
rect 1210 328 1266 362
rect 1300 328 1616 362
rect 1650 328 1706 362
rect 1740 328 1796 362
rect 1830 328 1886 362
rect 1920 328 1976 362
rect 2010 328 2066 362
rect 2100 328 2156 362
rect 2190 328 2246 362
rect 2280 328 2336 362
rect 2370 328 2426 362
rect 2460 328 2516 362
rect 2550 328 2606 362
rect 2640 328 2956 362
rect 2990 328 3046 362
rect 3080 328 3136 362
rect 3170 328 3226 362
rect 3260 328 3316 362
rect 3350 328 3406 362
rect 3440 328 3496 362
rect 3530 328 3586 362
rect 3620 328 3676 362
rect 3710 328 3766 362
rect 3800 328 3856 362
rect 3890 328 3946 362
rect 3980 328 4296 362
rect 4330 328 4386 362
rect 4420 328 4476 362
rect 4510 328 4566 362
rect 4600 328 4656 362
rect 4690 328 4746 362
rect 4780 328 4836 362
rect 4870 328 4926 362
rect 4960 328 5016 362
rect 5050 328 5106 362
rect 5140 328 5196 362
rect 5230 328 5286 362
rect 5320 328 5636 362
rect 5670 328 5726 362
rect 5760 328 5816 362
rect 5850 328 5906 362
rect 5940 328 5996 362
rect 6030 328 6086 362
rect 6120 328 6176 362
rect 6210 328 6266 362
rect 6300 328 6356 362
rect 6390 328 6446 362
rect 6480 328 6536 362
rect 6570 328 6626 362
rect 6660 328 6976 362
rect 7010 328 7066 362
rect 7100 328 7156 362
rect 7190 328 7246 362
rect 7280 328 7336 362
rect 7370 328 7426 362
rect 7460 328 7516 362
rect 7550 328 7606 362
rect 7640 328 7696 362
rect 7730 328 7786 362
rect 7820 328 7876 362
rect 7910 328 7966 362
rect 8000 328 8316 362
rect 8350 328 8406 362
rect 8440 328 8496 362
rect 8530 328 8586 362
rect 8620 328 8676 362
rect 8710 328 8766 362
rect 8800 328 8856 362
rect 8890 328 8946 362
rect 8980 328 9036 362
rect 9070 328 9126 362
rect 9160 328 9216 362
rect 9250 328 9306 362
rect 9340 328 9656 362
rect 9690 328 9746 362
rect 9780 328 9836 362
rect 9870 328 9926 362
rect 9960 328 10016 362
rect 10050 328 10106 362
rect 10140 328 10196 362
rect 10230 328 10286 362
rect 10320 328 10376 362
rect 10410 328 10466 362
rect 10500 328 10556 362
rect 10590 328 10646 362
rect 10680 328 10814 362
rect 146 296 10814 328
<< nsubdiff >>
rect 309 1402 1271 1421
rect 309 1368 440 1402
rect 474 1368 530 1402
rect 564 1368 620 1402
rect 654 1368 710 1402
rect 744 1368 800 1402
rect 834 1368 890 1402
rect 924 1368 980 1402
rect 1014 1368 1070 1402
rect 1104 1368 1160 1402
rect 1194 1368 1271 1402
rect 309 1349 1271 1368
rect 309 1345 381 1349
rect 309 1311 328 1345
rect 362 1311 381 1345
rect 309 1255 381 1311
rect 1199 1326 1271 1349
rect 1199 1292 1218 1326
rect 1252 1292 1271 1326
rect 309 1221 328 1255
rect 362 1221 381 1255
rect 309 1165 381 1221
rect 309 1131 328 1165
rect 362 1131 381 1165
rect 309 1075 381 1131
rect 309 1041 328 1075
rect 362 1041 381 1075
rect 309 985 381 1041
rect 309 951 328 985
rect 362 951 381 985
rect 309 895 381 951
rect 309 861 328 895
rect 362 861 381 895
rect 309 805 381 861
rect 309 771 328 805
rect 362 771 381 805
rect 309 715 381 771
rect 309 681 328 715
rect 362 681 381 715
rect 309 625 381 681
rect 309 591 328 625
rect 362 591 381 625
rect 1199 1236 1271 1292
rect 1199 1202 1218 1236
rect 1252 1202 1271 1236
rect 1199 1146 1271 1202
rect 1199 1112 1218 1146
rect 1252 1112 1271 1146
rect 1199 1056 1271 1112
rect 1199 1022 1218 1056
rect 1252 1022 1271 1056
rect 1199 966 1271 1022
rect 1199 932 1218 966
rect 1252 932 1271 966
rect 1199 876 1271 932
rect 1199 842 1218 876
rect 1252 842 1271 876
rect 1199 786 1271 842
rect 1199 752 1218 786
rect 1252 752 1271 786
rect 1199 696 1271 752
rect 1199 662 1218 696
rect 1252 662 1271 696
rect 1199 606 1271 662
rect 309 531 381 591
rect 1199 572 1218 606
rect 1252 572 1271 606
rect 1199 531 1271 572
rect 309 512 1271 531
rect 309 478 406 512
rect 440 478 496 512
rect 530 478 586 512
rect 620 478 676 512
rect 710 478 766 512
rect 800 478 856 512
rect 890 478 946 512
rect 980 478 1036 512
rect 1070 478 1126 512
rect 1160 478 1271 512
rect 309 459 1271 478
rect 1649 1402 2611 1421
rect 1649 1368 1780 1402
rect 1814 1368 1870 1402
rect 1904 1368 1960 1402
rect 1994 1368 2050 1402
rect 2084 1368 2140 1402
rect 2174 1368 2230 1402
rect 2264 1368 2320 1402
rect 2354 1368 2410 1402
rect 2444 1368 2500 1402
rect 2534 1368 2611 1402
rect 1649 1349 2611 1368
rect 1649 1345 1721 1349
rect 1649 1311 1668 1345
rect 1702 1311 1721 1345
rect 1649 1255 1721 1311
rect 2539 1326 2611 1349
rect 2539 1292 2558 1326
rect 2592 1292 2611 1326
rect 1649 1221 1668 1255
rect 1702 1221 1721 1255
rect 1649 1165 1721 1221
rect 1649 1131 1668 1165
rect 1702 1131 1721 1165
rect 1649 1075 1721 1131
rect 1649 1041 1668 1075
rect 1702 1041 1721 1075
rect 1649 985 1721 1041
rect 1649 951 1668 985
rect 1702 951 1721 985
rect 1649 895 1721 951
rect 1649 861 1668 895
rect 1702 861 1721 895
rect 1649 805 1721 861
rect 1649 771 1668 805
rect 1702 771 1721 805
rect 1649 715 1721 771
rect 1649 681 1668 715
rect 1702 681 1721 715
rect 1649 625 1721 681
rect 1649 591 1668 625
rect 1702 591 1721 625
rect 2539 1236 2611 1292
rect 2539 1202 2558 1236
rect 2592 1202 2611 1236
rect 2539 1146 2611 1202
rect 2539 1112 2558 1146
rect 2592 1112 2611 1146
rect 2539 1056 2611 1112
rect 2539 1022 2558 1056
rect 2592 1022 2611 1056
rect 2539 966 2611 1022
rect 2539 932 2558 966
rect 2592 932 2611 966
rect 2539 876 2611 932
rect 2539 842 2558 876
rect 2592 842 2611 876
rect 2539 786 2611 842
rect 2539 752 2558 786
rect 2592 752 2611 786
rect 2539 696 2611 752
rect 2539 662 2558 696
rect 2592 662 2611 696
rect 2539 606 2611 662
rect 1649 531 1721 591
rect 2539 572 2558 606
rect 2592 572 2611 606
rect 2539 531 2611 572
rect 1649 512 2611 531
rect 1649 478 1746 512
rect 1780 478 1836 512
rect 1870 478 1926 512
rect 1960 478 2016 512
rect 2050 478 2106 512
rect 2140 478 2196 512
rect 2230 478 2286 512
rect 2320 478 2376 512
rect 2410 478 2466 512
rect 2500 478 2611 512
rect 1649 459 2611 478
rect 2989 1402 3951 1421
rect 2989 1368 3120 1402
rect 3154 1368 3210 1402
rect 3244 1368 3300 1402
rect 3334 1368 3390 1402
rect 3424 1368 3480 1402
rect 3514 1368 3570 1402
rect 3604 1368 3660 1402
rect 3694 1368 3750 1402
rect 3784 1368 3840 1402
rect 3874 1368 3951 1402
rect 2989 1349 3951 1368
rect 2989 1345 3061 1349
rect 2989 1311 3008 1345
rect 3042 1311 3061 1345
rect 2989 1255 3061 1311
rect 3879 1326 3951 1349
rect 3879 1292 3898 1326
rect 3932 1292 3951 1326
rect 2989 1221 3008 1255
rect 3042 1221 3061 1255
rect 2989 1165 3061 1221
rect 2989 1131 3008 1165
rect 3042 1131 3061 1165
rect 2989 1075 3061 1131
rect 2989 1041 3008 1075
rect 3042 1041 3061 1075
rect 2989 985 3061 1041
rect 2989 951 3008 985
rect 3042 951 3061 985
rect 2989 895 3061 951
rect 2989 861 3008 895
rect 3042 861 3061 895
rect 2989 805 3061 861
rect 2989 771 3008 805
rect 3042 771 3061 805
rect 2989 715 3061 771
rect 2989 681 3008 715
rect 3042 681 3061 715
rect 2989 625 3061 681
rect 2989 591 3008 625
rect 3042 591 3061 625
rect 3879 1236 3951 1292
rect 3879 1202 3898 1236
rect 3932 1202 3951 1236
rect 3879 1146 3951 1202
rect 3879 1112 3898 1146
rect 3932 1112 3951 1146
rect 3879 1056 3951 1112
rect 3879 1022 3898 1056
rect 3932 1022 3951 1056
rect 3879 966 3951 1022
rect 3879 932 3898 966
rect 3932 932 3951 966
rect 3879 876 3951 932
rect 3879 842 3898 876
rect 3932 842 3951 876
rect 3879 786 3951 842
rect 3879 752 3898 786
rect 3932 752 3951 786
rect 3879 696 3951 752
rect 3879 662 3898 696
rect 3932 662 3951 696
rect 3879 606 3951 662
rect 2989 531 3061 591
rect 3879 572 3898 606
rect 3932 572 3951 606
rect 3879 531 3951 572
rect 2989 512 3951 531
rect 2989 478 3086 512
rect 3120 478 3176 512
rect 3210 478 3266 512
rect 3300 478 3356 512
rect 3390 478 3446 512
rect 3480 478 3536 512
rect 3570 478 3626 512
rect 3660 478 3716 512
rect 3750 478 3806 512
rect 3840 478 3951 512
rect 2989 459 3951 478
rect 4329 1402 5291 1421
rect 4329 1368 4460 1402
rect 4494 1368 4550 1402
rect 4584 1368 4640 1402
rect 4674 1368 4730 1402
rect 4764 1368 4820 1402
rect 4854 1368 4910 1402
rect 4944 1368 5000 1402
rect 5034 1368 5090 1402
rect 5124 1368 5180 1402
rect 5214 1368 5291 1402
rect 4329 1349 5291 1368
rect 4329 1345 4401 1349
rect 4329 1311 4348 1345
rect 4382 1311 4401 1345
rect 4329 1255 4401 1311
rect 5219 1326 5291 1349
rect 5219 1292 5238 1326
rect 5272 1292 5291 1326
rect 4329 1221 4348 1255
rect 4382 1221 4401 1255
rect 4329 1165 4401 1221
rect 4329 1131 4348 1165
rect 4382 1131 4401 1165
rect 4329 1075 4401 1131
rect 4329 1041 4348 1075
rect 4382 1041 4401 1075
rect 4329 985 4401 1041
rect 4329 951 4348 985
rect 4382 951 4401 985
rect 4329 895 4401 951
rect 4329 861 4348 895
rect 4382 861 4401 895
rect 4329 805 4401 861
rect 4329 771 4348 805
rect 4382 771 4401 805
rect 4329 715 4401 771
rect 4329 681 4348 715
rect 4382 681 4401 715
rect 4329 625 4401 681
rect 4329 591 4348 625
rect 4382 591 4401 625
rect 5219 1236 5291 1292
rect 5219 1202 5238 1236
rect 5272 1202 5291 1236
rect 5219 1146 5291 1202
rect 5219 1112 5238 1146
rect 5272 1112 5291 1146
rect 5219 1056 5291 1112
rect 5219 1022 5238 1056
rect 5272 1022 5291 1056
rect 5219 966 5291 1022
rect 5219 932 5238 966
rect 5272 932 5291 966
rect 5219 876 5291 932
rect 5219 842 5238 876
rect 5272 842 5291 876
rect 5219 786 5291 842
rect 5219 752 5238 786
rect 5272 752 5291 786
rect 5219 696 5291 752
rect 5219 662 5238 696
rect 5272 662 5291 696
rect 5219 606 5291 662
rect 4329 531 4401 591
rect 5219 572 5238 606
rect 5272 572 5291 606
rect 5219 531 5291 572
rect 4329 512 5291 531
rect 4329 478 4426 512
rect 4460 478 4516 512
rect 4550 478 4606 512
rect 4640 478 4696 512
rect 4730 478 4786 512
rect 4820 478 4876 512
rect 4910 478 4966 512
rect 5000 478 5056 512
rect 5090 478 5146 512
rect 5180 478 5291 512
rect 4329 459 5291 478
rect 5669 1402 6631 1421
rect 5669 1368 5800 1402
rect 5834 1368 5890 1402
rect 5924 1368 5980 1402
rect 6014 1368 6070 1402
rect 6104 1368 6160 1402
rect 6194 1368 6250 1402
rect 6284 1368 6340 1402
rect 6374 1368 6430 1402
rect 6464 1368 6520 1402
rect 6554 1368 6631 1402
rect 5669 1349 6631 1368
rect 5669 1345 5741 1349
rect 5669 1311 5688 1345
rect 5722 1311 5741 1345
rect 5669 1255 5741 1311
rect 6559 1326 6631 1349
rect 6559 1292 6578 1326
rect 6612 1292 6631 1326
rect 5669 1221 5688 1255
rect 5722 1221 5741 1255
rect 5669 1165 5741 1221
rect 5669 1131 5688 1165
rect 5722 1131 5741 1165
rect 5669 1075 5741 1131
rect 5669 1041 5688 1075
rect 5722 1041 5741 1075
rect 5669 985 5741 1041
rect 5669 951 5688 985
rect 5722 951 5741 985
rect 5669 895 5741 951
rect 5669 861 5688 895
rect 5722 861 5741 895
rect 5669 805 5741 861
rect 5669 771 5688 805
rect 5722 771 5741 805
rect 5669 715 5741 771
rect 5669 681 5688 715
rect 5722 681 5741 715
rect 5669 625 5741 681
rect 5669 591 5688 625
rect 5722 591 5741 625
rect 6559 1236 6631 1292
rect 6559 1202 6578 1236
rect 6612 1202 6631 1236
rect 6559 1146 6631 1202
rect 6559 1112 6578 1146
rect 6612 1112 6631 1146
rect 6559 1056 6631 1112
rect 6559 1022 6578 1056
rect 6612 1022 6631 1056
rect 6559 966 6631 1022
rect 6559 932 6578 966
rect 6612 932 6631 966
rect 6559 876 6631 932
rect 6559 842 6578 876
rect 6612 842 6631 876
rect 6559 786 6631 842
rect 6559 752 6578 786
rect 6612 752 6631 786
rect 6559 696 6631 752
rect 6559 662 6578 696
rect 6612 662 6631 696
rect 6559 606 6631 662
rect 5669 531 5741 591
rect 6559 572 6578 606
rect 6612 572 6631 606
rect 6559 531 6631 572
rect 5669 512 6631 531
rect 5669 478 5766 512
rect 5800 478 5856 512
rect 5890 478 5946 512
rect 5980 478 6036 512
rect 6070 478 6126 512
rect 6160 478 6216 512
rect 6250 478 6306 512
rect 6340 478 6396 512
rect 6430 478 6486 512
rect 6520 478 6631 512
rect 5669 459 6631 478
rect 7009 1402 7971 1421
rect 7009 1368 7140 1402
rect 7174 1368 7230 1402
rect 7264 1368 7320 1402
rect 7354 1368 7410 1402
rect 7444 1368 7500 1402
rect 7534 1368 7590 1402
rect 7624 1368 7680 1402
rect 7714 1368 7770 1402
rect 7804 1368 7860 1402
rect 7894 1368 7971 1402
rect 7009 1349 7971 1368
rect 7009 1345 7081 1349
rect 7009 1311 7028 1345
rect 7062 1311 7081 1345
rect 7009 1255 7081 1311
rect 7899 1326 7971 1349
rect 7899 1292 7918 1326
rect 7952 1292 7971 1326
rect 7009 1221 7028 1255
rect 7062 1221 7081 1255
rect 7009 1165 7081 1221
rect 7009 1131 7028 1165
rect 7062 1131 7081 1165
rect 7009 1075 7081 1131
rect 7009 1041 7028 1075
rect 7062 1041 7081 1075
rect 7009 985 7081 1041
rect 7009 951 7028 985
rect 7062 951 7081 985
rect 7009 895 7081 951
rect 7009 861 7028 895
rect 7062 861 7081 895
rect 7009 805 7081 861
rect 7009 771 7028 805
rect 7062 771 7081 805
rect 7009 715 7081 771
rect 7009 681 7028 715
rect 7062 681 7081 715
rect 7009 625 7081 681
rect 7009 591 7028 625
rect 7062 591 7081 625
rect 7899 1236 7971 1292
rect 7899 1202 7918 1236
rect 7952 1202 7971 1236
rect 7899 1146 7971 1202
rect 7899 1112 7918 1146
rect 7952 1112 7971 1146
rect 7899 1056 7971 1112
rect 7899 1022 7918 1056
rect 7952 1022 7971 1056
rect 7899 966 7971 1022
rect 7899 932 7918 966
rect 7952 932 7971 966
rect 7899 876 7971 932
rect 7899 842 7918 876
rect 7952 842 7971 876
rect 7899 786 7971 842
rect 7899 752 7918 786
rect 7952 752 7971 786
rect 7899 696 7971 752
rect 7899 662 7918 696
rect 7952 662 7971 696
rect 7899 606 7971 662
rect 7009 531 7081 591
rect 7899 572 7918 606
rect 7952 572 7971 606
rect 7899 531 7971 572
rect 7009 512 7971 531
rect 7009 478 7106 512
rect 7140 478 7196 512
rect 7230 478 7286 512
rect 7320 478 7376 512
rect 7410 478 7466 512
rect 7500 478 7556 512
rect 7590 478 7646 512
rect 7680 478 7736 512
rect 7770 478 7826 512
rect 7860 478 7971 512
rect 7009 459 7971 478
rect 8349 1402 9311 1421
rect 8349 1368 8480 1402
rect 8514 1368 8570 1402
rect 8604 1368 8660 1402
rect 8694 1368 8750 1402
rect 8784 1368 8840 1402
rect 8874 1368 8930 1402
rect 8964 1368 9020 1402
rect 9054 1368 9110 1402
rect 9144 1368 9200 1402
rect 9234 1368 9311 1402
rect 8349 1349 9311 1368
rect 8349 1345 8421 1349
rect 8349 1311 8368 1345
rect 8402 1311 8421 1345
rect 8349 1255 8421 1311
rect 9239 1326 9311 1349
rect 9239 1292 9258 1326
rect 9292 1292 9311 1326
rect 8349 1221 8368 1255
rect 8402 1221 8421 1255
rect 8349 1165 8421 1221
rect 8349 1131 8368 1165
rect 8402 1131 8421 1165
rect 8349 1075 8421 1131
rect 8349 1041 8368 1075
rect 8402 1041 8421 1075
rect 8349 985 8421 1041
rect 8349 951 8368 985
rect 8402 951 8421 985
rect 8349 895 8421 951
rect 8349 861 8368 895
rect 8402 861 8421 895
rect 8349 805 8421 861
rect 8349 771 8368 805
rect 8402 771 8421 805
rect 8349 715 8421 771
rect 8349 681 8368 715
rect 8402 681 8421 715
rect 8349 625 8421 681
rect 8349 591 8368 625
rect 8402 591 8421 625
rect 9239 1236 9311 1292
rect 9239 1202 9258 1236
rect 9292 1202 9311 1236
rect 9239 1146 9311 1202
rect 9239 1112 9258 1146
rect 9292 1112 9311 1146
rect 9239 1056 9311 1112
rect 9239 1022 9258 1056
rect 9292 1022 9311 1056
rect 9239 966 9311 1022
rect 9239 932 9258 966
rect 9292 932 9311 966
rect 9239 876 9311 932
rect 9239 842 9258 876
rect 9292 842 9311 876
rect 9239 786 9311 842
rect 9239 752 9258 786
rect 9292 752 9311 786
rect 9239 696 9311 752
rect 9239 662 9258 696
rect 9292 662 9311 696
rect 9239 606 9311 662
rect 8349 531 8421 591
rect 9239 572 9258 606
rect 9292 572 9311 606
rect 9239 531 9311 572
rect 8349 512 9311 531
rect 8349 478 8446 512
rect 8480 478 8536 512
rect 8570 478 8626 512
rect 8660 478 8716 512
rect 8750 478 8806 512
rect 8840 478 8896 512
rect 8930 478 8986 512
rect 9020 478 9076 512
rect 9110 478 9166 512
rect 9200 478 9311 512
rect 8349 459 9311 478
rect 9689 1402 10651 1421
rect 9689 1368 9820 1402
rect 9854 1368 9910 1402
rect 9944 1368 10000 1402
rect 10034 1368 10090 1402
rect 10124 1368 10180 1402
rect 10214 1368 10270 1402
rect 10304 1368 10360 1402
rect 10394 1368 10450 1402
rect 10484 1368 10540 1402
rect 10574 1368 10651 1402
rect 9689 1349 10651 1368
rect 9689 1345 9761 1349
rect 9689 1311 9708 1345
rect 9742 1311 9761 1345
rect 9689 1255 9761 1311
rect 10579 1326 10651 1349
rect 10579 1292 10598 1326
rect 10632 1292 10651 1326
rect 9689 1221 9708 1255
rect 9742 1221 9761 1255
rect 9689 1165 9761 1221
rect 9689 1131 9708 1165
rect 9742 1131 9761 1165
rect 9689 1075 9761 1131
rect 9689 1041 9708 1075
rect 9742 1041 9761 1075
rect 9689 985 9761 1041
rect 9689 951 9708 985
rect 9742 951 9761 985
rect 9689 895 9761 951
rect 9689 861 9708 895
rect 9742 861 9761 895
rect 9689 805 9761 861
rect 9689 771 9708 805
rect 9742 771 9761 805
rect 9689 715 9761 771
rect 9689 681 9708 715
rect 9742 681 9761 715
rect 9689 625 9761 681
rect 9689 591 9708 625
rect 9742 591 9761 625
rect 10579 1236 10651 1292
rect 10579 1202 10598 1236
rect 10632 1202 10651 1236
rect 10579 1146 10651 1202
rect 10579 1112 10598 1146
rect 10632 1112 10651 1146
rect 10579 1056 10651 1112
rect 10579 1022 10598 1056
rect 10632 1022 10651 1056
rect 10579 966 10651 1022
rect 10579 932 10598 966
rect 10632 932 10651 966
rect 10579 876 10651 932
rect 10579 842 10598 876
rect 10632 842 10651 876
rect 10579 786 10651 842
rect 10579 752 10598 786
rect 10632 752 10651 786
rect 10579 696 10651 752
rect 10579 662 10598 696
rect 10632 662 10651 696
rect 10579 606 10651 662
rect 9689 531 9761 591
rect 10579 572 10598 606
rect 10632 572 10651 606
rect 10579 531 10651 572
rect 9689 512 10651 531
rect 9689 478 9786 512
rect 9820 478 9876 512
rect 9910 478 9966 512
rect 10000 478 10056 512
rect 10090 478 10146 512
rect 10180 478 10236 512
rect 10270 478 10326 512
rect 10360 478 10416 512
rect 10450 478 10506 512
rect 10540 478 10651 512
rect 9689 459 10651 478
<< psubdiffcont >>
rect 180 1492 214 1526
rect 276 1515 310 1549
rect 366 1515 400 1549
rect 456 1515 490 1549
rect 546 1515 580 1549
rect 636 1515 670 1549
rect 726 1515 760 1549
rect 816 1515 850 1549
rect 906 1515 940 1549
rect 996 1515 1030 1549
rect 1086 1515 1120 1549
rect 1176 1515 1210 1549
rect 1266 1515 1300 1549
rect 1367 1492 1401 1526
rect 1520 1492 1554 1526
rect 1616 1515 1650 1549
rect 1706 1515 1740 1549
rect 1796 1515 1830 1549
rect 1886 1515 1920 1549
rect 1976 1515 2010 1549
rect 2066 1515 2100 1549
rect 2156 1515 2190 1549
rect 2246 1515 2280 1549
rect 2336 1515 2370 1549
rect 2426 1515 2460 1549
rect 2516 1515 2550 1549
rect 2606 1515 2640 1549
rect 2707 1492 2741 1526
rect 2860 1492 2894 1526
rect 2956 1515 2990 1549
rect 3046 1515 3080 1549
rect 3136 1515 3170 1549
rect 3226 1515 3260 1549
rect 3316 1515 3350 1549
rect 3406 1515 3440 1549
rect 3496 1515 3530 1549
rect 3586 1515 3620 1549
rect 3676 1515 3710 1549
rect 3766 1515 3800 1549
rect 3856 1515 3890 1549
rect 3946 1515 3980 1549
rect 4047 1492 4081 1526
rect 4200 1492 4234 1526
rect 4296 1515 4330 1549
rect 4386 1515 4420 1549
rect 4476 1515 4510 1549
rect 4566 1515 4600 1549
rect 4656 1515 4690 1549
rect 4746 1515 4780 1549
rect 4836 1515 4870 1549
rect 4926 1515 4960 1549
rect 5016 1515 5050 1549
rect 5106 1515 5140 1549
rect 5196 1515 5230 1549
rect 5286 1515 5320 1549
rect 5387 1492 5421 1526
rect 5540 1492 5574 1526
rect 5636 1515 5670 1549
rect 5726 1515 5760 1549
rect 5816 1515 5850 1549
rect 5906 1515 5940 1549
rect 5996 1515 6030 1549
rect 6086 1515 6120 1549
rect 6176 1515 6210 1549
rect 6266 1515 6300 1549
rect 6356 1515 6390 1549
rect 6446 1515 6480 1549
rect 6536 1515 6570 1549
rect 6626 1515 6660 1549
rect 6727 1492 6761 1526
rect 6880 1492 6914 1526
rect 6976 1515 7010 1549
rect 7066 1515 7100 1549
rect 7156 1515 7190 1549
rect 7246 1515 7280 1549
rect 7336 1515 7370 1549
rect 7426 1515 7460 1549
rect 7516 1515 7550 1549
rect 7606 1515 7640 1549
rect 7696 1515 7730 1549
rect 7786 1515 7820 1549
rect 7876 1515 7910 1549
rect 7966 1515 8000 1549
rect 8067 1492 8101 1526
rect 8220 1492 8254 1526
rect 8316 1515 8350 1549
rect 8406 1515 8440 1549
rect 8496 1515 8530 1549
rect 8586 1515 8620 1549
rect 8676 1515 8710 1549
rect 8766 1515 8800 1549
rect 8856 1515 8890 1549
rect 8946 1515 8980 1549
rect 9036 1515 9070 1549
rect 9126 1515 9160 1549
rect 9216 1515 9250 1549
rect 9306 1515 9340 1549
rect 9407 1492 9441 1526
rect 9560 1492 9594 1526
rect 9656 1515 9690 1549
rect 9746 1515 9780 1549
rect 9836 1515 9870 1549
rect 9926 1515 9960 1549
rect 10016 1515 10050 1549
rect 10106 1515 10140 1549
rect 10196 1515 10230 1549
rect 10286 1515 10320 1549
rect 10376 1515 10410 1549
rect 10466 1515 10500 1549
rect 10556 1515 10590 1549
rect 10646 1515 10680 1549
rect 10747 1492 10781 1526
rect 180 1402 214 1436
rect 180 1312 214 1346
rect 180 1222 214 1256
rect 180 1132 214 1166
rect 180 1042 214 1076
rect 180 952 214 986
rect 180 862 214 896
rect 180 772 214 806
rect 180 682 214 716
rect 180 592 214 626
rect 180 502 214 536
rect 1367 1402 1401 1436
rect 1520 1402 1554 1436
rect 1367 1312 1401 1346
rect 1520 1312 1554 1346
rect 1367 1222 1401 1256
rect 1520 1222 1554 1256
rect 1367 1132 1401 1166
rect 1520 1132 1554 1166
rect 1367 1042 1401 1076
rect 1520 1042 1554 1076
rect 1367 952 1401 986
rect 1520 952 1554 986
rect 1367 862 1401 896
rect 1520 862 1554 896
rect 1367 772 1401 806
rect 1520 772 1554 806
rect 1367 682 1401 716
rect 1520 682 1554 716
rect 1367 592 1401 626
rect 1520 592 1554 626
rect 1367 502 1401 536
rect 1520 502 1554 536
rect 180 412 214 446
rect 2707 1402 2741 1436
rect 2860 1402 2894 1436
rect 2707 1312 2741 1346
rect 2860 1312 2894 1346
rect 2707 1222 2741 1256
rect 2860 1222 2894 1256
rect 2707 1132 2741 1166
rect 2860 1132 2894 1166
rect 2707 1042 2741 1076
rect 2860 1042 2894 1076
rect 2707 952 2741 986
rect 2860 952 2894 986
rect 2707 862 2741 896
rect 2860 862 2894 896
rect 2707 772 2741 806
rect 2860 772 2894 806
rect 2707 682 2741 716
rect 2860 682 2894 716
rect 2707 592 2741 626
rect 2860 592 2894 626
rect 2707 502 2741 536
rect 2860 502 2894 536
rect 1367 412 1401 446
rect 1520 412 1554 446
rect 4047 1402 4081 1436
rect 4200 1402 4234 1436
rect 4047 1312 4081 1346
rect 4200 1312 4234 1346
rect 4047 1222 4081 1256
rect 4200 1222 4234 1256
rect 4047 1132 4081 1166
rect 4200 1132 4234 1166
rect 4047 1042 4081 1076
rect 4200 1042 4234 1076
rect 4047 952 4081 986
rect 4200 952 4234 986
rect 4047 862 4081 896
rect 4200 862 4234 896
rect 4047 772 4081 806
rect 4200 772 4234 806
rect 4047 682 4081 716
rect 4200 682 4234 716
rect 4047 592 4081 626
rect 4200 592 4234 626
rect 4047 502 4081 536
rect 4200 502 4234 536
rect 2707 412 2741 446
rect 2860 412 2894 446
rect 5387 1402 5421 1436
rect 5540 1402 5574 1436
rect 5387 1312 5421 1346
rect 5540 1312 5574 1346
rect 5387 1222 5421 1256
rect 5540 1222 5574 1256
rect 5387 1132 5421 1166
rect 5540 1132 5574 1166
rect 5387 1042 5421 1076
rect 5540 1042 5574 1076
rect 5387 952 5421 986
rect 5540 952 5574 986
rect 5387 862 5421 896
rect 5540 862 5574 896
rect 5387 772 5421 806
rect 5540 772 5574 806
rect 5387 682 5421 716
rect 5540 682 5574 716
rect 5387 592 5421 626
rect 5540 592 5574 626
rect 5387 502 5421 536
rect 5540 502 5574 536
rect 4047 412 4081 446
rect 4200 412 4234 446
rect 6727 1402 6761 1436
rect 6880 1402 6914 1436
rect 6727 1312 6761 1346
rect 6880 1312 6914 1346
rect 6727 1222 6761 1256
rect 6880 1222 6914 1256
rect 6727 1132 6761 1166
rect 6880 1132 6914 1166
rect 6727 1042 6761 1076
rect 6880 1042 6914 1076
rect 6727 952 6761 986
rect 6880 952 6914 986
rect 6727 862 6761 896
rect 6880 862 6914 896
rect 6727 772 6761 806
rect 6880 772 6914 806
rect 6727 682 6761 716
rect 6880 682 6914 716
rect 6727 592 6761 626
rect 6880 592 6914 626
rect 6727 502 6761 536
rect 6880 502 6914 536
rect 5387 412 5421 446
rect 5540 412 5574 446
rect 8067 1402 8101 1436
rect 8220 1402 8254 1436
rect 8067 1312 8101 1346
rect 8220 1312 8254 1346
rect 8067 1222 8101 1256
rect 8220 1222 8254 1256
rect 8067 1132 8101 1166
rect 8220 1132 8254 1166
rect 8067 1042 8101 1076
rect 8220 1042 8254 1076
rect 8067 952 8101 986
rect 8220 952 8254 986
rect 8067 862 8101 896
rect 8220 862 8254 896
rect 8067 772 8101 806
rect 8220 772 8254 806
rect 8067 682 8101 716
rect 8220 682 8254 716
rect 8067 592 8101 626
rect 8220 592 8254 626
rect 8067 502 8101 536
rect 8220 502 8254 536
rect 6727 412 6761 446
rect 6880 412 6914 446
rect 9407 1402 9441 1436
rect 9560 1402 9594 1436
rect 9407 1312 9441 1346
rect 9560 1312 9594 1346
rect 9407 1222 9441 1256
rect 9560 1222 9594 1256
rect 9407 1132 9441 1166
rect 9560 1132 9594 1166
rect 9407 1042 9441 1076
rect 9560 1042 9594 1076
rect 9407 952 9441 986
rect 9560 952 9594 986
rect 9407 862 9441 896
rect 9560 862 9594 896
rect 9407 772 9441 806
rect 9560 772 9594 806
rect 9407 682 9441 716
rect 9560 682 9594 716
rect 9407 592 9441 626
rect 9560 592 9594 626
rect 9407 502 9441 536
rect 9560 502 9594 536
rect 8067 412 8101 446
rect 8220 412 8254 446
rect 10747 1402 10781 1436
rect 10747 1312 10781 1346
rect 10747 1222 10781 1256
rect 10747 1132 10781 1166
rect 10747 1042 10781 1076
rect 10747 952 10781 986
rect 10747 862 10781 896
rect 10747 772 10781 806
rect 10747 682 10781 716
rect 10747 592 10781 626
rect 10747 502 10781 536
rect 9407 412 9441 446
rect 9560 412 9594 446
rect 10747 412 10781 446
rect 276 328 310 362
rect 366 328 400 362
rect 456 328 490 362
rect 546 328 580 362
rect 636 328 670 362
rect 726 328 760 362
rect 816 328 850 362
rect 906 328 940 362
rect 996 328 1030 362
rect 1086 328 1120 362
rect 1176 328 1210 362
rect 1266 328 1300 362
rect 1616 328 1650 362
rect 1706 328 1740 362
rect 1796 328 1830 362
rect 1886 328 1920 362
rect 1976 328 2010 362
rect 2066 328 2100 362
rect 2156 328 2190 362
rect 2246 328 2280 362
rect 2336 328 2370 362
rect 2426 328 2460 362
rect 2516 328 2550 362
rect 2606 328 2640 362
rect 2956 328 2990 362
rect 3046 328 3080 362
rect 3136 328 3170 362
rect 3226 328 3260 362
rect 3316 328 3350 362
rect 3406 328 3440 362
rect 3496 328 3530 362
rect 3586 328 3620 362
rect 3676 328 3710 362
rect 3766 328 3800 362
rect 3856 328 3890 362
rect 3946 328 3980 362
rect 4296 328 4330 362
rect 4386 328 4420 362
rect 4476 328 4510 362
rect 4566 328 4600 362
rect 4656 328 4690 362
rect 4746 328 4780 362
rect 4836 328 4870 362
rect 4926 328 4960 362
rect 5016 328 5050 362
rect 5106 328 5140 362
rect 5196 328 5230 362
rect 5286 328 5320 362
rect 5636 328 5670 362
rect 5726 328 5760 362
rect 5816 328 5850 362
rect 5906 328 5940 362
rect 5996 328 6030 362
rect 6086 328 6120 362
rect 6176 328 6210 362
rect 6266 328 6300 362
rect 6356 328 6390 362
rect 6446 328 6480 362
rect 6536 328 6570 362
rect 6626 328 6660 362
rect 6976 328 7010 362
rect 7066 328 7100 362
rect 7156 328 7190 362
rect 7246 328 7280 362
rect 7336 328 7370 362
rect 7426 328 7460 362
rect 7516 328 7550 362
rect 7606 328 7640 362
rect 7696 328 7730 362
rect 7786 328 7820 362
rect 7876 328 7910 362
rect 7966 328 8000 362
rect 8316 328 8350 362
rect 8406 328 8440 362
rect 8496 328 8530 362
rect 8586 328 8620 362
rect 8676 328 8710 362
rect 8766 328 8800 362
rect 8856 328 8890 362
rect 8946 328 8980 362
rect 9036 328 9070 362
rect 9126 328 9160 362
rect 9216 328 9250 362
rect 9306 328 9340 362
rect 9656 328 9690 362
rect 9746 328 9780 362
rect 9836 328 9870 362
rect 9926 328 9960 362
rect 10016 328 10050 362
rect 10106 328 10140 362
rect 10196 328 10230 362
rect 10286 328 10320 362
rect 10376 328 10410 362
rect 10466 328 10500 362
rect 10556 328 10590 362
rect 10646 328 10680 362
<< nsubdiffcont >>
rect 440 1368 474 1402
rect 530 1368 564 1402
rect 620 1368 654 1402
rect 710 1368 744 1402
rect 800 1368 834 1402
rect 890 1368 924 1402
rect 980 1368 1014 1402
rect 1070 1368 1104 1402
rect 1160 1368 1194 1402
rect 328 1311 362 1345
rect 1218 1292 1252 1326
rect 328 1221 362 1255
rect 328 1131 362 1165
rect 328 1041 362 1075
rect 328 951 362 985
rect 328 861 362 895
rect 328 771 362 805
rect 328 681 362 715
rect 328 591 362 625
rect 1218 1202 1252 1236
rect 1218 1112 1252 1146
rect 1218 1022 1252 1056
rect 1218 932 1252 966
rect 1218 842 1252 876
rect 1218 752 1252 786
rect 1218 662 1252 696
rect 1218 572 1252 606
rect 406 478 440 512
rect 496 478 530 512
rect 586 478 620 512
rect 676 478 710 512
rect 766 478 800 512
rect 856 478 890 512
rect 946 478 980 512
rect 1036 478 1070 512
rect 1126 478 1160 512
rect 1780 1368 1814 1402
rect 1870 1368 1904 1402
rect 1960 1368 1994 1402
rect 2050 1368 2084 1402
rect 2140 1368 2174 1402
rect 2230 1368 2264 1402
rect 2320 1368 2354 1402
rect 2410 1368 2444 1402
rect 2500 1368 2534 1402
rect 1668 1311 1702 1345
rect 2558 1292 2592 1326
rect 1668 1221 1702 1255
rect 1668 1131 1702 1165
rect 1668 1041 1702 1075
rect 1668 951 1702 985
rect 1668 861 1702 895
rect 1668 771 1702 805
rect 1668 681 1702 715
rect 1668 591 1702 625
rect 2558 1202 2592 1236
rect 2558 1112 2592 1146
rect 2558 1022 2592 1056
rect 2558 932 2592 966
rect 2558 842 2592 876
rect 2558 752 2592 786
rect 2558 662 2592 696
rect 2558 572 2592 606
rect 1746 478 1780 512
rect 1836 478 1870 512
rect 1926 478 1960 512
rect 2016 478 2050 512
rect 2106 478 2140 512
rect 2196 478 2230 512
rect 2286 478 2320 512
rect 2376 478 2410 512
rect 2466 478 2500 512
rect 3120 1368 3154 1402
rect 3210 1368 3244 1402
rect 3300 1368 3334 1402
rect 3390 1368 3424 1402
rect 3480 1368 3514 1402
rect 3570 1368 3604 1402
rect 3660 1368 3694 1402
rect 3750 1368 3784 1402
rect 3840 1368 3874 1402
rect 3008 1311 3042 1345
rect 3898 1292 3932 1326
rect 3008 1221 3042 1255
rect 3008 1131 3042 1165
rect 3008 1041 3042 1075
rect 3008 951 3042 985
rect 3008 861 3042 895
rect 3008 771 3042 805
rect 3008 681 3042 715
rect 3008 591 3042 625
rect 3898 1202 3932 1236
rect 3898 1112 3932 1146
rect 3898 1022 3932 1056
rect 3898 932 3932 966
rect 3898 842 3932 876
rect 3898 752 3932 786
rect 3898 662 3932 696
rect 3898 572 3932 606
rect 3086 478 3120 512
rect 3176 478 3210 512
rect 3266 478 3300 512
rect 3356 478 3390 512
rect 3446 478 3480 512
rect 3536 478 3570 512
rect 3626 478 3660 512
rect 3716 478 3750 512
rect 3806 478 3840 512
rect 4460 1368 4494 1402
rect 4550 1368 4584 1402
rect 4640 1368 4674 1402
rect 4730 1368 4764 1402
rect 4820 1368 4854 1402
rect 4910 1368 4944 1402
rect 5000 1368 5034 1402
rect 5090 1368 5124 1402
rect 5180 1368 5214 1402
rect 4348 1311 4382 1345
rect 5238 1292 5272 1326
rect 4348 1221 4382 1255
rect 4348 1131 4382 1165
rect 4348 1041 4382 1075
rect 4348 951 4382 985
rect 4348 861 4382 895
rect 4348 771 4382 805
rect 4348 681 4382 715
rect 4348 591 4382 625
rect 5238 1202 5272 1236
rect 5238 1112 5272 1146
rect 5238 1022 5272 1056
rect 5238 932 5272 966
rect 5238 842 5272 876
rect 5238 752 5272 786
rect 5238 662 5272 696
rect 5238 572 5272 606
rect 4426 478 4460 512
rect 4516 478 4550 512
rect 4606 478 4640 512
rect 4696 478 4730 512
rect 4786 478 4820 512
rect 4876 478 4910 512
rect 4966 478 5000 512
rect 5056 478 5090 512
rect 5146 478 5180 512
rect 5800 1368 5834 1402
rect 5890 1368 5924 1402
rect 5980 1368 6014 1402
rect 6070 1368 6104 1402
rect 6160 1368 6194 1402
rect 6250 1368 6284 1402
rect 6340 1368 6374 1402
rect 6430 1368 6464 1402
rect 6520 1368 6554 1402
rect 5688 1311 5722 1345
rect 6578 1292 6612 1326
rect 5688 1221 5722 1255
rect 5688 1131 5722 1165
rect 5688 1041 5722 1075
rect 5688 951 5722 985
rect 5688 861 5722 895
rect 5688 771 5722 805
rect 5688 681 5722 715
rect 5688 591 5722 625
rect 6578 1202 6612 1236
rect 6578 1112 6612 1146
rect 6578 1022 6612 1056
rect 6578 932 6612 966
rect 6578 842 6612 876
rect 6578 752 6612 786
rect 6578 662 6612 696
rect 6578 572 6612 606
rect 5766 478 5800 512
rect 5856 478 5890 512
rect 5946 478 5980 512
rect 6036 478 6070 512
rect 6126 478 6160 512
rect 6216 478 6250 512
rect 6306 478 6340 512
rect 6396 478 6430 512
rect 6486 478 6520 512
rect 7140 1368 7174 1402
rect 7230 1368 7264 1402
rect 7320 1368 7354 1402
rect 7410 1368 7444 1402
rect 7500 1368 7534 1402
rect 7590 1368 7624 1402
rect 7680 1368 7714 1402
rect 7770 1368 7804 1402
rect 7860 1368 7894 1402
rect 7028 1311 7062 1345
rect 7918 1292 7952 1326
rect 7028 1221 7062 1255
rect 7028 1131 7062 1165
rect 7028 1041 7062 1075
rect 7028 951 7062 985
rect 7028 861 7062 895
rect 7028 771 7062 805
rect 7028 681 7062 715
rect 7028 591 7062 625
rect 7918 1202 7952 1236
rect 7918 1112 7952 1146
rect 7918 1022 7952 1056
rect 7918 932 7952 966
rect 7918 842 7952 876
rect 7918 752 7952 786
rect 7918 662 7952 696
rect 7918 572 7952 606
rect 7106 478 7140 512
rect 7196 478 7230 512
rect 7286 478 7320 512
rect 7376 478 7410 512
rect 7466 478 7500 512
rect 7556 478 7590 512
rect 7646 478 7680 512
rect 7736 478 7770 512
rect 7826 478 7860 512
rect 8480 1368 8514 1402
rect 8570 1368 8604 1402
rect 8660 1368 8694 1402
rect 8750 1368 8784 1402
rect 8840 1368 8874 1402
rect 8930 1368 8964 1402
rect 9020 1368 9054 1402
rect 9110 1368 9144 1402
rect 9200 1368 9234 1402
rect 8368 1311 8402 1345
rect 9258 1292 9292 1326
rect 8368 1221 8402 1255
rect 8368 1131 8402 1165
rect 8368 1041 8402 1075
rect 8368 951 8402 985
rect 8368 861 8402 895
rect 8368 771 8402 805
rect 8368 681 8402 715
rect 8368 591 8402 625
rect 9258 1202 9292 1236
rect 9258 1112 9292 1146
rect 9258 1022 9292 1056
rect 9258 932 9292 966
rect 9258 842 9292 876
rect 9258 752 9292 786
rect 9258 662 9292 696
rect 9258 572 9292 606
rect 8446 478 8480 512
rect 8536 478 8570 512
rect 8626 478 8660 512
rect 8716 478 8750 512
rect 8806 478 8840 512
rect 8896 478 8930 512
rect 8986 478 9020 512
rect 9076 478 9110 512
rect 9166 478 9200 512
rect 9820 1368 9854 1402
rect 9910 1368 9944 1402
rect 10000 1368 10034 1402
rect 10090 1368 10124 1402
rect 10180 1368 10214 1402
rect 10270 1368 10304 1402
rect 10360 1368 10394 1402
rect 10450 1368 10484 1402
rect 10540 1368 10574 1402
rect 9708 1311 9742 1345
rect 10598 1292 10632 1326
rect 9708 1221 9742 1255
rect 9708 1131 9742 1165
rect 9708 1041 9742 1075
rect 9708 951 9742 985
rect 9708 861 9742 895
rect 9708 771 9742 805
rect 9708 681 9742 715
rect 9708 591 9742 625
rect 10598 1202 10632 1236
rect 10598 1112 10632 1146
rect 10598 1022 10632 1056
rect 10598 932 10632 966
rect 10598 842 10632 876
rect 10598 752 10632 786
rect 10598 662 10632 696
rect 10598 572 10632 606
rect 9786 478 9820 512
rect 9876 478 9910 512
rect 9966 478 10000 512
rect 10056 478 10090 512
rect 10146 478 10180 512
rect 10236 478 10270 512
rect 10326 478 10360 512
rect 10416 478 10450 512
rect 10506 478 10540 512
<< locali >>
rect 120 1897 10840 1910
rect 120 1863 303 1897
rect 337 1863 503 1897
rect 537 1863 703 1897
rect 737 1863 903 1897
rect 937 1863 1103 1897
rect 1137 1863 1303 1897
rect 1337 1863 1503 1897
rect 1537 1863 1703 1897
rect 1737 1863 1903 1897
rect 1937 1863 2103 1897
rect 2137 1863 2303 1897
rect 2337 1863 2503 1897
rect 2537 1863 2703 1897
rect 2737 1863 2903 1897
rect 2937 1863 3103 1897
rect 3137 1863 3303 1897
rect 3337 1863 3503 1897
rect 3537 1863 3703 1897
rect 3737 1863 3903 1897
rect 3937 1863 4103 1897
rect 4137 1863 4303 1897
rect 4337 1863 4503 1897
rect 4537 1863 4703 1897
rect 4737 1863 4903 1897
rect 4937 1863 5103 1897
rect 5137 1863 5303 1897
rect 5337 1863 5503 1897
rect 5537 1863 5703 1897
rect 5737 1863 5903 1897
rect 5937 1863 6103 1897
rect 6137 1863 6303 1897
rect 6337 1863 6503 1897
rect 6537 1863 6703 1897
rect 6737 1863 6903 1897
rect 6937 1863 7103 1897
rect 7137 1863 7303 1897
rect 7337 1863 7503 1897
rect 7537 1863 7703 1897
rect 7737 1863 7903 1897
rect 7937 1863 8103 1897
rect 8137 1863 8303 1897
rect 8337 1863 8503 1897
rect 8537 1863 8703 1897
rect 8737 1863 8903 1897
rect 8937 1863 9103 1897
rect 9137 1863 9303 1897
rect 9337 1863 9503 1897
rect 9537 1863 9703 1897
rect 9737 1863 9903 1897
rect 9937 1863 10103 1897
rect 10137 1863 10303 1897
rect 10337 1863 10503 1897
rect 10537 1863 10703 1897
rect 10737 1863 10840 1897
rect 120 1850 10840 1863
rect 146 1564 10814 1584
rect 146 1530 166 1564
rect 200 1530 256 1564
rect 290 1549 346 1564
rect 380 1549 436 1564
rect 470 1549 526 1564
rect 560 1549 616 1564
rect 650 1549 706 1564
rect 740 1549 796 1564
rect 830 1549 886 1564
rect 920 1549 976 1564
rect 1010 1549 1066 1564
rect 1100 1549 1156 1564
rect 1190 1549 1246 1564
rect 1280 1549 1336 1564
rect 310 1530 346 1549
rect 400 1530 436 1549
rect 490 1530 526 1549
rect 580 1530 616 1549
rect 670 1530 706 1549
rect 760 1530 796 1549
rect 850 1530 886 1549
rect 940 1530 976 1549
rect 1030 1530 1066 1549
rect 1120 1530 1156 1549
rect 1210 1530 1246 1549
rect 1300 1530 1336 1549
rect 1370 1530 1506 1564
rect 1540 1530 1596 1564
rect 1630 1549 1686 1564
rect 1720 1549 1776 1564
rect 1810 1549 1866 1564
rect 1900 1549 1956 1564
rect 1990 1549 2046 1564
rect 2080 1549 2136 1564
rect 2170 1549 2226 1564
rect 2260 1549 2316 1564
rect 2350 1549 2406 1564
rect 2440 1549 2496 1564
rect 2530 1549 2586 1564
rect 2620 1549 2676 1564
rect 1650 1530 1686 1549
rect 1740 1530 1776 1549
rect 1830 1530 1866 1549
rect 1920 1530 1956 1549
rect 2010 1530 2046 1549
rect 2100 1530 2136 1549
rect 2190 1530 2226 1549
rect 2280 1530 2316 1549
rect 2370 1530 2406 1549
rect 2460 1530 2496 1549
rect 2550 1530 2586 1549
rect 2640 1530 2676 1549
rect 2710 1530 2846 1564
rect 2880 1530 2936 1564
rect 2970 1549 3026 1564
rect 3060 1549 3116 1564
rect 3150 1549 3206 1564
rect 3240 1549 3296 1564
rect 3330 1549 3386 1564
rect 3420 1549 3476 1564
rect 3510 1549 3566 1564
rect 3600 1549 3656 1564
rect 3690 1549 3746 1564
rect 3780 1549 3836 1564
rect 3870 1549 3926 1564
rect 3960 1549 4016 1564
rect 2990 1530 3026 1549
rect 3080 1530 3116 1549
rect 3170 1530 3206 1549
rect 3260 1530 3296 1549
rect 3350 1530 3386 1549
rect 3440 1530 3476 1549
rect 3530 1530 3566 1549
rect 3620 1530 3656 1549
rect 3710 1530 3746 1549
rect 3800 1530 3836 1549
rect 3890 1530 3926 1549
rect 3980 1530 4016 1549
rect 4050 1530 4186 1564
rect 4220 1530 4276 1564
rect 4310 1549 4366 1564
rect 4400 1549 4456 1564
rect 4490 1549 4546 1564
rect 4580 1549 4636 1564
rect 4670 1549 4726 1564
rect 4760 1549 4816 1564
rect 4850 1549 4906 1564
rect 4940 1549 4996 1564
rect 5030 1549 5086 1564
rect 5120 1549 5176 1564
rect 5210 1549 5266 1564
rect 5300 1549 5356 1564
rect 4330 1530 4366 1549
rect 4420 1530 4456 1549
rect 4510 1530 4546 1549
rect 4600 1530 4636 1549
rect 4690 1530 4726 1549
rect 4780 1530 4816 1549
rect 4870 1530 4906 1549
rect 4960 1530 4996 1549
rect 5050 1530 5086 1549
rect 5140 1530 5176 1549
rect 5230 1530 5266 1549
rect 5320 1530 5356 1549
rect 5390 1530 5526 1564
rect 5560 1530 5616 1564
rect 5650 1549 5706 1564
rect 5740 1549 5796 1564
rect 5830 1549 5886 1564
rect 5920 1549 5976 1564
rect 6010 1549 6066 1564
rect 6100 1549 6156 1564
rect 6190 1549 6246 1564
rect 6280 1549 6336 1564
rect 6370 1549 6426 1564
rect 6460 1549 6516 1564
rect 6550 1549 6606 1564
rect 6640 1549 6696 1564
rect 5670 1530 5706 1549
rect 5760 1530 5796 1549
rect 5850 1530 5886 1549
rect 5940 1530 5976 1549
rect 6030 1530 6066 1549
rect 6120 1530 6156 1549
rect 6210 1530 6246 1549
rect 6300 1530 6336 1549
rect 6390 1530 6426 1549
rect 6480 1530 6516 1549
rect 6570 1530 6606 1549
rect 6660 1530 6696 1549
rect 6730 1530 6866 1564
rect 6900 1530 6956 1564
rect 6990 1549 7046 1564
rect 7080 1549 7136 1564
rect 7170 1549 7226 1564
rect 7260 1549 7316 1564
rect 7350 1549 7406 1564
rect 7440 1549 7496 1564
rect 7530 1549 7586 1564
rect 7620 1549 7676 1564
rect 7710 1549 7766 1564
rect 7800 1549 7856 1564
rect 7890 1549 7946 1564
rect 7980 1549 8036 1564
rect 7010 1530 7046 1549
rect 7100 1530 7136 1549
rect 7190 1530 7226 1549
rect 7280 1530 7316 1549
rect 7370 1530 7406 1549
rect 7460 1530 7496 1549
rect 7550 1530 7586 1549
rect 7640 1530 7676 1549
rect 7730 1530 7766 1549
rect 7820 1530 7856 1549
rect 7910 1530 7946 1549
rect 8000 1530 8036 1549
rect 8070 1530 8206 1564
rect 8240 1530 8296 1564
rect 8330 1549 8386 1564
rect 8420 1549 8476 1564
rect 8510 1549 8566 1564
rect 8600 1549 8656 1564
rect 8690 1549 8746 1564
rect 8780 1549 8836 1564
rect 8870 1549 8926 1564
rect 8960 1549 9016 1564
rect 9050 1549 9106 1564
rect 9140 1549 9196 1564
rect 9230 1549 9286 1564
rect 9320 1549 9376 1564
rect 8350 1530 8386 1549
rect 8440 1530 8476 1549
rect 8530 1530 8566 1549
rect 8620 1530 8656 1549
rect 8710 1530 8746 1549
rect 8800 1530 8836 1549
rect 8890 1530 8926 1549
rect 8980 1530 9016 1549
rect 9070 1530 9106 1549
rect 9160 1530 9196 1549
rect 9250 1530 9286 1549
rect 9340 1530 9376 1549
rect 9410 1530 9546 1564
rect 9580 1530 9636 1564
rect 9670 1549 9726 1564
rect 9760 1549 9816 1564
rect 9850 1549 9906 1564
rect 9940 1549 9996 1564
rect 10030 1549 10086 1564
rect 10120 1549 10176 1564
rect 10210 1549 10266 1564
rect 10300 1549 10356 1564
rect 10390 1549 10446 1564
rect 10480 1549 10536 1564
rect 10570 1549 10626 1564
rect 10660 1549 10716 1564
rect 9690 1530 9726 1549
rect 9780 1530 9816 1549
rect 9870 1530 9906 1549
rect 9960 1530 9996 1549
rect 10050 1530 10086 1549
rect 10140 1530 10176 1549
rect 10230 1530 10266 1549
rect 10320 1530 10356 1549
rect 10410 1530 10446 1549
rect 10500 1530 10536 1549
rect 10590 1530 10626 1549
rect 10680 1530 10716 1549
rect 10750 1530 10814 1564
rect 146 1526 276 1530
rect 146 1492 180 1526
rect 214 1515 276 1526
rect 310 1515 366 1530
rect 400 1515 456 1530
rect 490 1515 546 1530
rect 580 1515 636 1530
rect 670 1515 726 1530
rect 760 1515 816 1530
rect 850 1515 906 1530
rect 940 1515 996 1530
rect 1030 1515 1086 1530
rect 1120 1515 1176 1530
rect 1210 1515 1266 1530
rect 1300 1526 1616 1530
rect 1300 1515 1367 1526
rect 214 1492 1367 1515
rect 1401 1492 1520 1526
rect 1554 1515 1616 1526
rect 1650 1515 1706 1530
rect 1740 1515 1796 1530
rect 1830 1515 1886 1530
rect 1920 1515 1976 1530
rect 2010 1515 2066 1530
rect 2100 1515 2156 1530
rect 2190 1515 2246 1530
rect 2280 1515 2336 1530
rect 2370 1515 2426 1530
rect 2460 1515 2516 1530
rect 2550 1515 2606 1530
rect 2640 1526 2956 1530
rect 2640 1515 2707 1526
rect 1554 1492 2707 1515
rect 2741 1492 2860 1526
rect 2894 1515 2956 1526
rect 2990 1515 3046 1530
rect 3080 1515 3136 1530
rect 3170 1515 3226 1530
rect 3260 1515 3316 1530
rect 3350 1515 3406 1530
rect 3440 1515 3496 1530
rect 3530 1515 3586 1530
rect 3620 1515 3676 1530
rect 3710 1515 3766 1530
rect 3800 1515 3856 1530
rect 3890 1515 3946 1530
rect 3980 1526 4296 1530
rect 3980 1515 4047 1526
rect 2894 1492 4047 1515
rect 4081 1492 4200 1526
rect 4234 1515 4296 1526
rect 4330 1515 4386 1530
rect 4420 1515 4476 1530
rect 4510 1515 4566 1530
rect 4600 1515 4656 1530
rect 4690 1515 4746 1530
rect 4780 1515 4836 1530
rect 4870 1515 4926 1530
rect 4960 1515 5016 1530
rect 5050 1515 5106 1530
rect 5140 1515 5196 1530
rect 5230 1515 5286 1530
rect 5320 1526 5636 1530
rect 5320 1515 5387 1526
rect 4234 1492 5387 1515
rect 5421 1492 5540 1526
rect 5574 1515 5636 1526
rect 5670 1515 5726 1530
rect 5760 1515 5816 1530
rect 5850 1515 5906 1530
rect 5940 1515 5996 1530
rect 6030 1515 6086 1530
rect 6120 1515 6176 1530
rect 6210 1515 6266 1530
rect 6300 1515 6356 1530
rect 6390 1515 6446 1530
rect 6480 1515 6536 1530
rect 6570 1515 6626 1530
rect 6660 1526 6976 1530
rect 6660 1515 6727 1526
rect 5574 1492 6727 1515
rect 6761 1492 6880 1526
rect 6914 1515 6976 1526
rect 7010 1515 7066 1530
rect 7100 1515 7156 1530
rect 7190 1515 7246 1530
rect 7280 1515 7336 1530
rect 7370 1515 7426 1530
rect 7460 1515 7516 1530
rect 7550 1515 7606 1530
rect 7640 1515 7696 1530
rect 7730 1515 7786 1530
rect 7820 1515 7876 1530
rect 7910 1515 7966 1530
rect 8000 1526 8316 1530
rect 8000 1515 8067 1526
rect 6914 1492 8067 1515
rect 8101 1492 8220 1526
rect 8254 1515 8316 1526
rect 8350 1515 8406 1530
rect 8440 1515 8496 1530
rect 8530 1515 8586 1530
rect 8620 1515 8676 1530
rect 8710 1515 8766 1530
rect 8800 1515 8856 1530
rect 8890 1515 8946 1530
rect 8980 1515 9036 1530
rect 9070 1515 9126 1530
rect 9160 1515 9216 1530
rect 9250 1515 9306 1530
rect 9340 1526 9656 1530
rect 9340 1515 9407 1526
rect 8254 1492 9407 1515
rect 9441 1492 9560 1526
rect 9594 1515 9656 1526
rect 9690 1515 9746 1530
rect 9780 1515 9836 1530
rect 9870 1515 9926 1530
rect 9960 1515 10016 1530
rect 10050 1515 10106 1530
rect 10140 1515 10196 1530
rect 10230 1515 10286 1530
rect 10320 1515 10376 1530
rect 10410 1515 10466 1530
rect 10500 1515 10556 1530
rect 10590 1515 10646 1530
rect 10680 1526 10814 1530
rect 10680 1515 10747 1526
rect 9594 1492 10747 1515
rect 10781 1492 10814 1526
rect 146 1485 10814 1492
rect 146 1436 245 1485
rect 146 1402 180 1436
rect 214 1402 245 1436
rect 1335 1436 1585 1485
rect 146 1346 245 1402
rect 146 1312 180 1346
rect 214 1312 245 1346
rect 146 1256 245 1312
rect 146 1222 180 1256
rect 214 1222 245 1256
rect 146 1166 245 1222
rect 146 1132 180 1166
rect 214 1132 245 1166
rect 146 1076 245 1132
rect 146 1042 180 1076
rect 214 1042 245 1076
rect 146 986 245 1042
rect 146 952 180 986
rect 214 952 245 986
rect 146 896 245 952
rect 146 862 180 896
rect 214 862 245 896
rect 146 806 245 862
rect 146 772 180 806
rect 214 772 245 806
rect 146 716 245 772
rect 146 682 180 716
rect 214 682 245 716
rect 146 626 245 682
rect 146 592 180 626
rect 214 592 245 626
rect 146 536 245 592
rect 146 502 180 536
rect 214 502 245 536
rect 146 446 245 502
rect 309 1404 1271 1421
rect 309 1370 330 1404
rect 364 1370 420 1404
rect 454 1402 510 1404
rect 544 1402 600 1404
rect 634 1402 690 1404
rect 724 1402 780 1404
rect 814 1402 870 1404
rect 904 1402 960 1404
rect 994 1402 1050 1404
rect 1084 1402 1140 1404
rect 1174 1402 1230 1404
rect 474 1370 510 1402
rect 564 1370 600 1402
rect 654 1370 690 1402
rect 744 1370 780 1402
rect 834 1370 870 1402
rect 924 1370 960 1402
rect 1014 1370 1050 1402
rect 1104 1370 1140 1402
rect 1194 1370 1230 1402
rect 1264 1370 1271 1404
rect 309 1368 440 1370
rect 474 1368 530 1370
rect 564 1368 620 1370
rect 654 1368 710 1370
rect 744 1368 800 1370
rect 834 1368 890 1370
rect 924 1368 980 1370
rect 1014 1368 1070 1370
rect 1104 1368 1160 1370
rect 1194 1368 1271 1370
rect 309 1349 1271 1368
rect 309 1345 381 1349
rect 309 1311 328 1345
rect 362 1311 381 1345
rect 309 1255 381 1311
rect 1199 1326 1271 1349
rect 1199 1292 1218 1326
rect 1252 1292 1271 1326
rect 309 1221 328 1255
rect 362 1221 381 1255
rect 309 1165 381 1221
rect 309 1131 328 1165
rect 362 1131 381 1165
rect 309 1075 381 1131
rect 309 1041 328 1075
rect 362 1041 381 1075
rect 309 985 381 1041
rect 309 951 328 985
rect 362 951 381 985
rect 309 895 381 951
rect 309 861 328 895
rect 362 861 381 895
rect 309 805 381 861
rect 309 771 328 805
rect 362 771 381 805
rect 309 715 381 771
rect 309 681 328 715
rect 362 681 381 715
rect 309 625 381 681
rect 309 591 328 625
rect 362 591 381 625
rect 443 1228 1137 1287
rect 443 1194 504 1228
rect 538 1200 594 1228
rect 628 1200 684 1228
rect 718 1200 774 1228
rect 550 1194 594 1200
rect 650 1194 684 1200
rect 750 1194 774 1200
rect 808 1200 864 1228
rect 808 1194 816 1200
rect 443 1166 516 1194
rect 550 1166 616 1194
rect 650 1166 716 1194
rect 750 1166 816 1194
rect 850 1194 864 1200
rect 898 1200 954 1228
rect 898 1194 916 1200
rect 850 1166 916 1194
rect 950 1194 954 1200
rect 988 1200 1044 1228
rect 988 1194 1016 1200
rect 1078 1194 1137 1228
rect 950 1166 1016 1194
rect 1050 1166 1137 1194
rect 443 1138 1137 1166
rect 443 1104 504 1138
rect 538 1104 594 1138
rect 628 1104 684 1138
rect 718 1104 774 1138
rect 808 1104 864 1138
rect 898 1104 954 1138
rect 988 1104 1044 1138
rect 1078 1104 1137 1138
rect 443 1100 1137 1104
rect 443 1066 516 1100
rect 550 1066 616 1100
rect 650 1066 716 1100
rect 750 1066 816 1100
rect 850 1066 916 1100
rect 950 1066 1016 1100
rect 1050 1066 1137 1100
rect 443 1048 1137 1066
rect 443 1014 504 1048
rect 538 1014 594 1048
rect 628 1014 684 1048
rect 718 1014 774 1048
rect 808 1014 864 1048
rect 898 1014 954 1048
rect 988 1014 1044 1048
rect 1078 1014 1137 1048
rect 443 1000 1137 1014
rect 443 966 516 1000
rect 550 966 616 1000
rect 650 966 716 1000
rect 750 966 816 1000
rect 850 966 916 1000
rect 950 966 1016 1000
rect 1050 966 1137 1000
rect 443 958 1137 966
rect 443 924 504 958
rect 538 924 594 958
rect 628 924 684 958
rect 718 924 774 958
rect 808 924 864 958
rect 898 924 954 958
rect 988 924 1044 958
rect 1078 924 1137 958
rect 443 900 1137 924
rect 443 868 516 900
rect 550 868 616 900
rect 650 868 716 900
rect 750 868 816 900
rect 443 834 504 868
rect 550 866 594 868
rect 650 866 684 868
rect 750 866 774 868
rect 538 834 594 866
rect 628 834 684 866
rect 718 834 774 866
rect 808 866 816 868
rect 850 868 916 900
rect 850 866 864 868
rect 808 834 864 866
rect 898 866 916 868
rect 950 868 1016 900
rect 1050 868 1137 900
rect 950 866 954 868
rect 898 834 954 866
rect 988 866 1016 868
rect 988 834 1044 866
rect 1078 834 1137 868
rect 443 800 1137 834
rect 443 778 516 800
rect 550 778 616 800
rect 650 778 716 800
rect 750 778 816 800
rect 443 744 504 778
rect 550 766 594 778
rect 650 766 684 778
rect 750 766 774 778
rect 538 744 594 766
rect 628 744 684 766
rect 718 744 774 766
rect 808 766 816 778
rect 850 778 916 800
rect 850 766 864 778
rect 808 744 864 766
rect 898 766 916 778
rect 950 778 1016 800
rect 1050 778 1137 800
rect 950 766 954 778
rect 898 744 954 766
rect 988 766 1016 778
rect 988 744 1044 766
rect 1078 744 1137 778
rect 443 700 1137 744
rect 443 688 516 700
rect 550 688 616 700
rect 650 688 716 700
rect 750 688 816 700
rect 443 654 504 688
rect 550 666 594 688
rect 650 666 684 688
rect 750 666 774 688
rect 538 654 594 666
rect 628 654 684 666
rect 718 654 774 666
rect 808 666 816 688
rect 850 688 916 700
rect 850 666 864 688
rect 808 654 864 666
rect 898 666 916 688
rect 950 688 1016 700
rect 1050 688 1137 700
rect 950 666 954 688
rect 898 654 954 666
rect 988 666 1016 688
rect 988 654 1044 666
rect 1078 654 1137 688
rect 443 593 1137 654
rect 1199 1236 1271 1292
rect 1199 1202 1218 1236
rect 1252 1202 1271 1236
rect 1199 1146 1271 1202
rect 1199 1112 1218 1146
rect 1252 1112 1271 1146
rect 1199 1056 1271 1112
rect 1199 1022 1218 1056
rect 1252 1022 1271 1056
rect 1199 966 1271 1022
rect 1199 932 1218 966
rect 1252 932 1271 966
rect 1199 876 1271 932
rect 1199 842 1218 876
rect 1252 842 1271 876
rect 1199 786 1271 842
rect 1199 752 1218 786
rect 1252 752 1271 786
rect 1199 696 1271 752
rect 1199 662 1218 696
rect 1252 662 1271 696
rect 1199 606 1271 662
rect 309 531 381 591
rect 1199 572 1218 606
rect 1252 572 1271 606
rect 1199 531 1271 572
rect 309 512 1271 531
rect 309 478 406 512
rect 440 478 496 512
rect 530 478 586 512
rect 620 478 676 512
rect 710 478 766 512
rect 800 478 856 512
rect 890 478 946 512
rect 980 478 1036 512
rect 1070 478 1126 512
rect 1160 478 1271 512
rect 309 459 1271 478
rect 1335 1402 1367 1436
rect 1401 1402 1520 1436
rect 1554 1402 1585 1436
rect 2675 1436 2925 1485
rect 1335 1346 1585 1402
rect 1335 1312 1367 1346
rect 1401 1312 1520 1346
rect 1554 1312 1585 1346
rect 1335 1256 1585 1312
rect 1335 1222 1367 1256
rect 1401 1222 1520 1256
rect 1554 1222 1585 1256
rect 1335 1166 1585 1222
rect 1335 1132 1367 1166
rect 1401 1132 1520 1166
rect 1554 1132 1585 1166
rect 1335 1076 1585 1132
rect 1335 1042 1367 1076
rect 1401 1042 1520 1076
rect 1554 1042 1585 1076
rect 1335 986 1585 1042
rect 1335 952 1367 986
rect 1401 952 1520 986
rect 1554 952 1585 986
rect 1335 896 1585 952
rect 1335 862 1367 896
rect 1401 862 1520 896
rect 1554 862 1585 896
rect 1335 806 1585 862
rect 1335 772 1367 806
rect 1401 772 1520 806
rect 1554 772 1585 806
rect 1335 716 1585 772
rect 1335 682 1367 716
rect 1401 682 1520 716
rect 1554 682 1585 716
rect 1335 626 1585 682
rect 1335 592 1367 626
rect 1401 592 1520 626
rect 1554 592 1585 626
rect 1335 536 1585 592
rect 1335 502 1367 536
rect 1401 502 1520 536
rect 1554 502 1585 536
rect 146 412 180 446
rect 214 412 245 446
rect 146 395 245 412
rect 1335 446 1585 502
rect 1649 1404 2611 1421
rect 1649 1370 1670 1404
rect 1704 1370 1760 1404
rect 1794 1402 1850 1404
rect 1884 1402 1940 1404
rect 1974 1402 2030 1404
rect 2064 1402 2120 1404
rect 2154 1402 2210 1404
rect 2244 1402 2300 1404
rect 2334 1402 2390 1404
rect 2424 1402 2480 1404
rect 2514 1402 2570 1404
rect 1814 1370 1850 1402
rect 1904 1370 1940 1402
rect 1994 1370 2030 1402
rect 2084 1370 2120 1402
rect 2174 1370 2210 1402
rect 2264 1370 2300 1402
rect 2354 1370 2390 1402
rect 2444 1370 2480 1402
rect 2534 1370 2570 1402
rect 2604 1370 2611 1404
rect 1649 1368 1780 1370
rect 1814 1368 1870 1370
rect 1904 1368 1960 1370
rect 1994 1368 2050 1370
rect 2084 1368 2140 1370
rect 2174 1368 2230 1370
rect 2264 1368 2320 1370
rect 2354 1368 2410 1370
rect 2444 1368 2500 1370
rect 2534 1368 2611 1370
rect 1649 1349 2611 1368
rect 1649 1345 1721 1349
rect 1649 1311 1668 1345
rect 1702 1311 1721 1345
rect 1649 1255 1721 1311
rect 2539 1326 2611 1349
rect 2539 1292 2558 1326
rect 2592 1292 2611 1326
rect 1649 1221 1668 1255
rect 1702 1221 1721 1255
rect 1649 1165 1721 1221
rect 1649 1131 1668 1165
rect 1702 1131 1721 1165
rect 1649 1075 1721 1131
rect 1649 1041 1668 1075
rect 1702 1041 1721 1075
rect 1649 985 1721 1041
rect 1649 951 1668 985
rect 1702 951 1721 985
rect 1649 895 1721 951
rect 1649 861 1668 895
rect 1702 861 1721 895
rect 1649 805 1721 861
rect 1649 771 1668 805
rect 1702 771 1721 805
rect 1649 715 1721 771
rect 1649 681 1668 715
rect 1702 681 1721 715
rect 1649 625 1721 681
rect 1649 591 1668 625
rect 1702 591 1721 625
rect 1783 1228 2477 1287
rect 1783 1194 1844 1228
rect 1878 1200 1934 1228
rect 1968 1200 2024 1228
rect 2058 1200 2114 1228
rect 1890 1194 1934 1200
rect 1990 1194 2024 1200
rect 2090 1194 2114 1200
rect 2148 1200 2204 1228
rect 2148 1194 2156 1200
rect 1783 1166 1856 1194
rect 1890 1166 1956 1194
rect 1990 1166 2056 1194
rect 2090 1166 2156 1194
rect 2190 1194 2204 1200
rect 2238 1200 2294 1228
rect 2238 1194 2256 1200
rect 2190 1166 2256 1194
rect 2290 1194 2294 1200
rect 2328 1200 2384 1228
rect 2328 1194 2356 1200
rect 2418 1194 2477 1228
rect 2290 1166 2356 1194
rect 2390 1166 2477 1194
rect 1783 1138 2477 1166
rect 1783 1104 1844 1138
rect 1878 1104 1934 1138
rect 1968 1104 2024 1138
rect 2058 1104 2114 1138
rect 2148 1104 2204 1138
rect 2238 1104 2294 1138
rect 2328 1104 2384 1138
rect 2418 1104 2477 1138
rect 1783 1100 2477 1104
rect 1783 1066 1856 1100
rect 1890 1066 1956 1100
rect 1990 1066 2056 1100
rect 2090 1066 2156 1100
rect 2190 1066 2256 1100
rect 2290 1066 2356 1100
rect 2390 1066 2477 1100
rect 1783 1048 2477 1066
rect 1783 1014 1844 1048
rect 1878 1014 1934 1048
rect 1968 1014 2024 1048
rect 2058 1014 2114 1048
rect 2148 1014 2204 1048
rect 2238 1014 2294 1048
rect 2328 1014 2384 1048
rect 2418 1014 2477 1048
rect 1783 1000 2477 1014
rect 1783 966 1856 1000
rect 1890 966 1956 1000
rect 1990 966 2056 1000
rect 2090 966 2156 1000
rect 2190 966 2256 1000
rect 2290 966 2356 1000
rect 2390 966 2477 1000
rect 1783 958 2477 966
rect 1783 924 1844 958
rect 1878 924 1934 958
rect 1968 924 2024 958
rect 2058 924 2114 958
rect 2148 924 2204 958
rect 2238 924 2294 958
rect 2328 924 2384 958
rect 2418 924 2477 958
rect 1783 900 2477 924
rect 1783 868 1856 900
rect 1890 868 1956 900
rect 1990 868 2056 900
rect 2090 868 2156 900
rect 1783 834 1844 868
rect 1890 866 1934 868
rect 1990 866 2024 868
rect 2090 866 2114 868
rect 1878 834 1934 866
rect 1968 834 2024 866
rect 2058 834 2114 866
rect 2148 866 2156 868
rect 2190 868 2256 900
rect 2190 866 2204 868
rect 2148 834 2204 866
rect 2238 866 2256 868
rect 2290 868 2356 900
rect 2390 868 2477 900
rect 2290 866 2294 868
rect 2238 834 2294 866
rect 2328 866 2356 868
rect 2328 834 2384 866
rect 2418 834 2477 868
rect 1783 800 2477 834
rect 1783 778 1856 800
rect 1890 778 1956 800
rect 1990 778 2056 800
rect 2090 778 2156 800
rect 1783 744 1844 778
rect 1890 766 1934 778
rect 1990 766 2024 778
rect 2090 766 2114 778
rect 1878 744 1934 766
rect 1968 744 2024 766
rect 2058 744 2114 766
rect 2148 766 2156 778
rect 2190 778 2256 800
rect 2190 766 2204 778
rect 2148 744 2204 766
rect 2238 766 2256 778
rect 2290 778 2356 800
rect 2390 778 2477 800
rect 2290 766 2294 778
rect 2238 744 2294 766
rect 2328 766 2356 778
rect 2328 744 2384 766
rect 2418 744 2477 778
rect 1783 700 2477 744
rect 1783 688 1856 700
rect 1890 688 1956 700
rect 1990 688 2056 700
rect 2090 688 2156 700
rect 1783 654 1844 688
rect 1890 666 1934 688
rect 1990 666 2024 688
rect 2090 666 2114 688
rect 1878 654 1934 666
rect 1968 654 2024 666
rect 2058 654 2114 666
rect 2148 666 2156 688
rect 2190 688 2256 700
rect 2190 666 2204 688
rect 2148 654 2204 666
rect 2238 666 2256 688
rect 2290 688 2356 700
rect 2390 688 2477 700
rect 2290 666 2294 688
rect 2238 654 2294 666
rect 2328 666 2356 688
rect 2328 654 2384 666
rect 2418 654 2477 688
rect 1783 593 2477 654
rect 2539 1236 2611 1292
rect 2539 1202 2558 1236
rect 2592 1202 2611 1236
rect 2539 1146 2611 1202
rect 2539 1112 2558 1146
rect 2592 1112 2611 1146
rect 2539 1056 2611 1112
rect 2539 1022 2558 1056
rect 2592 1022 2611 1056
rect 2539 966 2611 1022
rect 2539 932 2558 966
rect 2592 932 2611 966
rect 2539 876 2611 932
rect 2539 842 2558 876
rect 2592 842 2611 876
rect 2539 786 2611 842
rect 2539 752 2558 786
rect 2592 752 2611 786
rect 2539 696 2611 752
rect 2539 662 2558 696
rect 2592 662 2611 696
rect 2539 606 2611 662
rect 1649 531 1721 591
rect 2539 572 2558 606
rect 2592 572 2611 606
rect 2539 531 2611 572
rect 1649 512 2611 531
rect 1649 478 1746 512
rect 1780 478 1836 512
rect 1870 478 1926 512
rect 1960 478 2016 512
rect 2050 478 2106 512
rect 2140 478 2196 512
rect 2230 478 2286 512
rect 2320 478 2376 512
rect 2410 478 2466 512
rect 2500 478 2611 512
rect 1649 459 2611 478
rect 2675 1402 2707 1436
rect 2741 1402 2860 1436
rect 2894 1402 2925 1436
rect 4015 1436 4265 1485
rect 2675 1346 2925 1402
rect 2675 1312 2707 1346
rect 2741 1312 2860 1346
rect 2894 1312 2925 1346
rect 2675 1256 2925 1312
rect 2675 1222 2707 1256
rect 2741 1222 2860 1256
rect 2894 1222 2925 1256
rect 2675 1166 2925 1222
rect 2675 1132 2707 1166
rect 2741 1132 2860 1166
rect 2894 1132 2925 1166
rect 2675 1076 2925 1132
rect 2675 1042 2707 1076
rect 2741 1042 2860 1076
rect 2894 1042 2925 1076
rect 2675 986 2925 1042
rect 2675 952 2707 986
rect 2741 952 2860 986
rect 2894 952 2925 986
rect 2675 896 2925 952
rect 2675 862 2707 896
rect 2741 862 2860 896
rect 2894 862 2925 896
rect 2675 806 2925 862
rect 2675 772 2707 806
rect 2741 772 2860 806
rect 2894 772 2925 806
rect 2675 716 2925 772
rect 2675 682 2707 716
rect 2741 682 2860 716
rect 2894 682 2925 716
rect 2675 626 2925 682
rect 2675 592 2707 626
rect 2741 592 2860 626
rect 2894 592 2925 626
rect 2675 536 2925 592
rect 2675 502 2707 536
rect 2741 502 2860 536
rect 2894 502 2925 536
rect 1335 412 1367 446
rect 1401 412 1520 446
rect 1554 412 1585 446
rect 1335 395 1585 412
rect 2675 446 2925 502
rect 2989 1404 3951 1421
rect 2989 1370 3010 1404
rect 3044 1370 3100 1404
rect 3134 1402 3190 1404
rect 3224 1402 3280 1404
rect 3314 1402 3370 1404
rect 3404 1402 3460 1404
rect 3494 1402 3550 1404
rect 3584 1402 3640 1404
rect 3674 1402 3730 1404
rect 3764 1402 3820 1404
rect 3854 1402 3910 1404
rect 3154 1370 3190 1402
rect 3244 1370 3280 1402
rect 3334 1370 3370 1402
rect 3424 1370 3460 1402
rect 3514 1370 3550 1402
rect 3604 1370 3640 1402
rect 3694 1370 3730 1402
rect 3784 1370 3820 1402
rect 3874 1370 3910 1402
rect 3944 1370 3951 1404
rect 2989 1368 3120 1370
rect 3154 1368 3210 1370
rect 3244 1368 3300 1370
rect 3334 1368 3390 1370
rect 3424 1368 3480 1370
rect 3514 1368 3570 1370
rect 3604 1368 3660 1370
rect 3694 1368 3750 1370
rect 3784 1368 3840 1370
rect 3874 1368 3951 1370
rect 2989 1349 3951 1368
rect 2989 1345 3061 1349
rect 2989 1311 3008 1345
rect 3042 1311 3061 1345
rect 2989 1255 3061 1311
rect 3879 1326 3951 1349
rect 3879 1292 3898 1326
rect 3932 1292 3951 1326
rect 2989 1221 3008 1255
rect 3042 1221 3061 1255
rect 2989 1165 3061 1221
rect 2989 1131 3008 1165
rect 3042 1131 3061 1165
rect 2989 1075 3061 1131
rect 2989 1041 3008 1075
rect 3042 1041 3061 1075
rect 2989 985 3061 1041
rect 2989 951 3008 985
rect 3042 951 3061 985
rect 2989 895 3061 951
rect 2989 861 3008 895
rect 3042 861 3061 895
rect 2989 805 3061 861
rect 2989 771 3008 805
rect 3042 771 3061 805
rect 2989 715 3061 771
rect 2989 681 3008 715
rect 3042 681 3061 715
rect 2989 625 3061 681
rect 2989 591 3008 625
rect 3042 591 3061 625
rect 3123 1228 3817 1287
rect 3123 1194 3184 1228
rect 3218 1200 3274 1228
rect 3308 1200 3364 1228
rect 3398 1200 3454 1228
rect 3230 1194 3274 1200
rect 3330 1194 3364 1200
rect 3430 1194 3454 1200
rect 3488 1200 3544 1228
rect 3488 1194 3496 1200
rect 3123 1166 3196 1194
rect 3230 1166 3296 1194
rect 3330 1166 3396 1194
rect 3430 1166 3496 1194
rect 3530 1194 3544 1200
rect 3578 1200 3634 1228
rect 3578 1194 3596 1200
rect 3530 1166 3596 1194
rect 3630 1194 3634 1200
rect 3668 1200 3724 1228
rect 3668 1194 3696 1200
rect 3758 1194 3817 1228
rect 3630 1166 3696 1194
rect 3730 1166 3817 1194
rect 3123 1138 3817 1166
rect 3123 1104 3184 1138
rect 3218 1104 3274 1138
rect 3308 1104 3364 1138
rect 3398 1104 3454 1138
rect 3488 1104 3544 1138
rect 3578 1104 3634 1138
rect 3668 1104 3724 1138
rect 3758 1104 3817 1138
rect 3123 1100 3817 1104
rect 3123 1066 3196 1100
rect 3230 1066 3296 1100
rect 3330 1066 3396 1100
rect 3430 1066 3496 1100
rect 3530 1066 3596 1100
rect 3630 1066 3696 1100
rect 3730 1066 3817 1100
rect 3123 1048 3817 1066
rect 3123 1014 3184 1048
rect 3218 1014 3274 1048
rect 3308 1014 3364 1048
rect 3398 1014 3454 1048
rect 3488 1014 3544 1048
rect 3578 1014 3634 1048
rect 3668 1014 3724 1048
rect 3758 1014 3817 1048
rect 3123 1000 3817 1014
rect 3123 966 3196 1000
rect 3230 966 3296 1000
rect 3330 966 3396 1000
rect 3430 966 3496 1000
rect 3530 966 3596 1000
rect 3630 966 3696 1000
rect 3730 966 3817 1000
rect 3123 958 3817 966
rect 3123 924 3184 958
rect 3218 924 3274 958
rect 3308 924 3364 958
rect 3398 924 3454 958
rect 3488 924 3544 958
rect 3578 924 3634 958
rect 3668 924 3724 958
rect 3758 924 3817 958
rect 3123 900 3817 924
rect 3123 868 3196 900
rect 3230 868 3296 900
rect 3330 868 3396 900
rect 3430 868 3496 900
rect 3123 834 3184 868
rect 3230 866 3274 868
rect 3330 866 3364 868
rect 3430 866 3454 868
rect 3218 834 3274 866
rect 3308 834 3364 866
rect 3398 834 3454 866
rect 3488 866 3496 868
rect 3530 868 3596 900
rect 3530 866 3544 868
rect 3488 834 3544 866
rect 3578 866 3596 868
rect 3630 868 3696 900
rect 3730 868 3817 900
rect 3630 866 3634 868
rect 3578 834 3634 866
rect 3668 866 3696 868
rect 3668 834 3724 866
rect 3758 834 3817 868
rect 3123 800 3817 834
rect 3123 778 3196 800
rect 3230 778 3296 800
rect 3330 778 3396 800
rect 3430 778 3496 800
rect 3123 744 3184 778
rect 3230 766 3274 778
rect 3330 766 3364 778
rect 3430 766 3454 778
rect 3218 744 3274 766
rect 3308 744 3364 766
rect 3398 744 3454 766
rect 3488 766 3496 778
rect 3530 778 3596 800
rect 3530 766 3544 778
rect 3488 744 3544 766
rect 3578 766 3596 778
rect 3630 778 3696 800
rect 3730 778 3817 800
rect 3630 766 3634 778
rect 3578 744 3634 766
rect 3668 766 3696 778
rect 3668 744 3724 766
rect 3758 744 3817 778
rect 3123 700 3817 744
rect 3123 688 3196 700
rect 3230 688 3296 700
rect 3330 688 3396 700
rect 3430 688 3496 700
rect 3123 654 3184 688
rect 3230 666 3274 688
rect 3330 666 3364 688
rect 3430 666 3454 688
rect 3218 654 3274 666
rect 3308 654 3364 666
rect 3398 654 3454 666
rect 3488 666 3496 688
rect 3530 688 3596 700
rect 3530 666 3544 688
rect 3488 654 3544 666
rect 3578 666 3596 688
rect 3630 688 3696 700
rect 3730 688 3817 700
rect 3630 666 3634 688
rect 3578 654 3634 666
rect 3668 666 3696 688
rect 3668 654 3724 666
rect 3758 654 3817 688
rect 3123 593 3817 654
rect 3879 1236 3951 1292
rect 3879 1202 3898 1236
rect 3932 1202 3951 1236
rect 3879 1146 3951 1202
rect 3879 1112 3898 1146
rect 3932 1112 3951 1146
rect 3879 1056 3951 1112
rect 3879 1022 3898 1056
rect 3932 1022 3951 1056
rect 3879 966 3951 1022
rect 3879 932 3898 966
rect 3932 932 3951 966
rect 3879 876 3951 932
rect 3879 842 3898 876
rect 3932 842 3951 876
rect 3879 786 3951 842
rect 3879 752 3898 786
rect 3932 752 3951 786
rect 3879 696 3951 752
rect 3879 662 3898 696
rect 3932 662 3951 696
rect 3879 606 3951 662
rect 2989 531 3061 591
rect 3879 572 3898 606
rect 3932 572 3951 606
rect 3879 531 3951 572
rect 2989 512 3951 531
rect 2989 478 3086 512
rect 3120 478 3176 512
rect 3210 478 3266 512
rect 3300 478 3356 512
rect 3390 478 3446 512
rect 3480 478 3536 512
rect 3570 478 3626 512
rect 3660 478 3716 512
rect 3750 478 3806 512
rect 3840 478 3951 512
rect 2989 459 3951 478
rect 4015 1402 4047 1436
rect 4081 1402 4200 1436
rect 4234 1402 4265 1436
rect 5355 1436 5605 1485
rect 4015 1346 4265 1402
rect 4015 1312 4047 1346
rect 4081 1312 4200 1346
rect 4234 1312 4265 1346
rect 4015 1256 4265 1312
rect 4015 1222 4047 1256
rect 4081 1222 4200 1256
rect 4234 1222 4265 1256
rect 4015 1166 4265 1222
rect 4015 1132 4047 1166
rect 4081 1132 4200 1166
rect 4234 1132 4265 1166
rect 4015 1076 4265 1132
rect 4015 1042 4047 1076
rect 4081 1042 4200 1076
rect 4234 1042 4265 1076
rect 4015 986 4265 1042
rect 4015 952 4047 986
rect 4081 952 4200 986
rect 4234 952 4265 986
rect 4015 896 4265 952
rect 4015 862 4047 896
rect 4081 862 4200 896
rect 4234 862 4265 896
rect 4015 806 4265 862
rect 4015 772 4047 806
rect 4081 772 4200 806
rect 4234 772 4265 806
rect 4015 716 4265 772
rect 4015 682 4047 716
rect 4081 682 4200 716
rect 4234 682 4265 716
rect 4015 626 4265 682
rect 4015 592 4047 626
rect 4081 592 4200 626
rect 4234 592 4265 626
rect 4015 536 4265 592
rect 4015 502 4047 536
rect 4081 502 4200 536
rect 4234 502 4265 536
rect 2675 412 2707 446
rect 2741 412 2860 446
rect 2894 412 2925 446
rect 2675 395 2925 412
rect 4015 446 4265 502
rect 4329 1404 5291 1421
rect 4329 1370 4350 1404
rect 4384 1370 4440 1404
rect 4474 1402 4530 1404
rect 4564 1402 4620 1404
rect 4654 1402 4710 1404
rect 4744 1402 4800 1404
rect 4834 1402 4890 1404
rect 4924 1402 4980 1404
rect 5014 1402 5070 1404
rect 5104 1402 5160 1404
rect 5194 1402 5250 1404
rect 4494 1370 4530 1402
rect 4584 1370 4620 1402
rect 4674 1370 4710 1402
rect 4764 1370 4800 1402
rect 4854 1370 4890 1402
rect 4944 1370 4980 1402
rect 5034 1370 5070 1402
rect 5124 1370 5160 1402
rect 5214 1370 5250 1402
rect 5284 1370 5291 1404
rect 4329 1368 4460 1370
rect 4494 1368 4550 1370
rect 4584 1368 4640 1370
rect 4674 1368 4730 1370
rect 4764 1368 4820 1370
rect 4854 1368 4910 1370
rect 4944 1368 5000 1370
rect 5034 1368 5090 1370
rect 5124 1368 5180 1370
rect 5214 1368 5291 1370
rect 4329 1349 5291 1368
rect 4329 1345 4401 1349
rect 4329 1311 4348 1345
rect 4382 1311 4401 1345
rect 4329 1255 4401 1311
rect 5219 1326 5291 1349
rect 5219 1292 5238 1326
rect 5272 1292 5291 1326
rect 4329 1221 4348 1255
rect 4382 1221 4401 1255
rect 4329 1165 4401 1221
rect 4329 1131 4348 1165
rect 4382 1131 4401 1165
rect 4329 1075 4401 1131
rect 4329 1041 4348 1075
rect 4382 1041 4401 1075
rect 4329 985 4401 1041
rect 4329 951 4348 985
rect 4382 951 4401 985
rect 4329 895 4401 951
rect 4329 861 4348 895
rect 4382 861 4401 895
rect 4329 805 4401 861
rect 4329 771 4348 805
rect 4382 771 4401 805
rect 4329 715 4401 771
rect 4329 681 4348 715
rect 4382 681 4401 715
rect 4329 625 4401 681
rect 4329 591 4348 625
rect 4382 591 4401 625
rect 4463 1228 5157 1287
rect 4463 1194 4524 1228
rect 4558 1200 4614 1228
rect 4648 1200 4704 1228
rect 4738 1200 4794 1228
rect 4570 1194 4614 1200
rect 4670 1194 4704 1200
rect 4770 1194 4794 1200
rect 4828 1200 4884 1228
rect 4828 1194 4836 1200
rect 4463 1166 4536 1194
rect 4570 1166 4636 1194
rect 4670 1166 4736 1194
rect 4770 1166 4836 1194
rect 4870 1194 4884 1200
rect 4918 1200 4974 1228
rect 4918 1194 4936 1200
rect 4870 1166 4936 1194
rect 4970 1194 4974 1200
rect 5008 1200 5064 1228
rect 5008 1194 5036 1200
rect 5098 1194 5157 1228
rect 4970 1166 5036 1194
rect 5070 1166 5157 1194
rect 4463 1138 5157 1166
rect 4463 1104 4524 1138
rect 4558 1104 4614 1138
rect 4648 1104 4704 1138
rect 4738 1104 4794 1138
rect 4828 1104 4884 1138
rect 4918 1104 4974 1138
rect 5008 1104 5064 1138
rect 5098 1104 5157 1138
rect 4463 1100 5157 1104
rect 4463 1066 4536 1100
rect 4570 1066 4636 1100
rect 4670 1066 4736 1100
rect 4770 1066 4836 1100
rect 4870 1066 4936 1100
rect 4970 1066 5036 1100
rect 5070 1066 5157 1100
rect 4463 1048 5157 1066
rect 4463 1014 4524 1048
rect 4558 1014 4614 1048
rect 4648 1014 4704 1048
rect 4738 1014 4794 1048
rect 4828 1014 4884 1048
rect 4918 1014 4974 1048
rect 5008 1014 5064 1048
rect 5098 1014 5157 1048
rect 4463 1000 5157 1014
rect 4463 966 4536 1000
rect 4570 966 4636 1000
rect 4670 966 4736 1000
rect 4770 966 4836 1000
rect 4870 966 4936 1000
rect 4970 966 5036 1000
rect 5070 966 5157 1000
rect 4463 958 5157 966
rect 4463 924 4524 958
rect 4558 924 4614 958
rect 4648 924 4704 958
rect 4738 924 4794 958
rect 4828 924 4884 958
rect 4918 924 4974 958
rect 5008 924 5064 958
rect 5098 924 5157 958
rect 4463 900 5157 924
rect 4463 868 4536 900
rect 4570 868 4636 900
rect 4670 868 4736 900
rect 4770 868 4836 900
rect 4463 834 4524 868
rect 4570 866 4614 868
rect 4670 866 4704 868
rect 4770 866 4794 868
rect 4558 834 4614 866
rect 4648 834 4704 866
rect 4738 834 4794 866
rect 4828 866 4836 868
rect 4870 868 4936 900
rect 4870 866 4884 868
rect 4828 834 4884 866
rect 4918 866 4936 868
rect 4970 868 5036 900
rect 5070 868 5157 900
rect 4970 866 4974 868
rect 4918 834 4974 866
rect 5008 866 5036 868
rect 5008 834 5064 866
rect 5098 834 5157 868
rect 4463 800 5157 834
rect 4463 778 4536 800
rect 4570 778 4636 800
rect 4670 778 4736 800
rect 4770 778 4836 800
rect 4463 744 4524 778
rect 4570 766 4614 778
rect 4670 766 4704 778
rect 4770 766 4794 778
rect 4558 744 4614 766
rect 4648 744 4704 766
rect 4738 744 4794 766
rect 4828 766 4836 778
rect 4870 778 4936 800
rect 4870 766 4884 778
rect 4828 744 4884 766
rect 4918 766 4936 778
rect 4970 778 5036 800
rect 5070 778 5157 800
rect 4970 766 4974 778
rect 4918 744 4974 766
rect 5008 766 5036 778
rect 5008 744 5064 766
rect 5098 744 5157 778
rect 4463 700 5157 744
rect 4463 688 4536 700
rect 4570 688 4636 700
rect 4670 688 4736 700
rect 4770 688 4836 700
rect 4463 654 4524 688
rect 4570 666 4614 688
rect 4670 666 4704 688
rect 4770 666 4794 688
rect 4558 654 4614 666
rect 4648 654 4704 666
rect 4738 654 4794 666
rect 4828 666 4836 688
rect 4870 688 4936 700
rect 4870 666 4884 688
rect 4828 654 4884 666
rect 4918 666 4936 688
rect 4970 688 5036 700
rect 5070 688 5157 700
rect 4970 666 4974 688
rect 4918 654 4974 666
rect 5008 666 5036 688
rect 5008 654 5064 666
rect 5098 654 5157 688
rect 4463 593 5157 654
rect 5219 1236 5291 1292
rect 5219 1202 5238 1236
rect 5272 1202 5291 1236
rect 5219 1146 5291 1202
rect 5219 1112 5238 1146
rect 5272 1112 5291 1146
rect 5219 1056 5291 1112
rect 5219 1022 5238 1056
rect 5272 1022 5291 1056
rect 5219 966 5291 1022
rect 5219 932 5238 966
rect 5272 932 5291 966
rect 5219 876 5291 932
rect 5219 842 5238 876
rect 5272 842 5291 876
rect 5219 786 5291 842
rect 5219 752 5238 786
rect 5272 752 5291 786
rect 5219 696 5291 752
rect 5219 662 5238 696
rect 5272 662 5291 696
rect 5219 606 5291 662
rect 4329 531 4401 591
rect 5219 572 5238 606
rect 5272 572 5291 606
rect 5219 531 5291 572
rect 4329 512 5291 531
rect 4329 478 4426 512
rect 4460 478 4516 512
rect 4550 478 4606 512
rect 4640 478 4696 512
rect 4730 478 4786 512
rect 4820 478 4876 512
rect 4910 478 4966 512
rect 5000 478 5056 512
rect 5090 478 5146 512
rect 5180 478 5291 512
rect 4329 459 5291 478
rect 5355 1402 5387 1436
rect 5421 1402 5540 1436
rect 5574 1402 5605 1436
rect 6695 1436 6945 1485
rect 5355 1346 5605 1402
rect 5355 1312 5387 1346
rect 5421 1312 5540 1346
rect 5574 1312 5605 1346
rect 5355 1256 5605 1312
rect 5355 1222 5387 1256
rect 5421 1222 5540 1256
rect 5574 1222 5605 1256
rect 5355 1166 5605 1222
rect 5355 1132 5387 1166
rect 5421 1132 5540 1166
rect 5574 1132 5605 1166
rect 5355 1076 5605 1132
rect 5355 1042 5387 1076
rect 5421 1042 5540 1076
rect 5574 1042 5605 1076
rect 5355 986 5605 1042
rect 5355 952 5387 986
rect 5421 952 5540 986
rect 5574 952 5605 986
rect 5355 896 5605 952
rect 5355 862 5387 896
rect 5421 862 5540 896
rect 5574 862 5605 896
rect 5355 806 5605 862
rect 5355 772 5387 806
rect 5421 772 5540 806
rect 5574 772 5605 806
rect 5355 716 5605 772
rect 5355 682 5387 716
rect 5421 682 5540 716
rect 5574 682 5605 716
rect 5355 626 5605 682
rect 5355 592 5387 626
rect 5421 592 5540 626
rect 5574 592 5605 626
rect 5355 536 5605 592
rect 5355 502 5387 536
rect 5421 502 5540 536
rect 5574 502 5605 536
rect 4015 412 4047 446
rect 4081 412 4200 446
rect 4234 412 4265 446
rect 4015 395 4265 412
rect 5355 446 5605 502
rect 5669 1404 6631 1421
rect 5669 1370 5690 1404
rect 5724 1370 5780 1404
rect 5814 1402 5870 1404
rect 5904 1402 5960 1404
rect 5994 1402 6050 1404
rect 6084 1402 6140 1404
rect 6174 1402 6230 1404
rect 6264 1402 6320 1404
rect 6354 1402 6410 1404
rect 6444 1402 6500 1404
rect 6534 1402 6590 1404
rect 5834 1370 5870 1402
rect 5924 1370 5960 1402
rect 6014 1370 6050 1402
rect 6104 1370 6140 1402
rect 6194 1370 6230 1402
rect 6284 1370 6320 1402
rect 6374 1370 6410 1402
rect 6464 1370 6500 1402
rect 6554 1370 6590 1402
rect 6624 1370 6631 1404
rect 5669 1368 5800 1370
rect 5834 1368 5890 1370
rect 5924 1368 5980 1370
rect 6014 1368 6070 1370
rect 6104 1368 6160 1370
rect 6194 1368 6250 1370
rect 6284 1368 6340 1370
rect 6374 1368 6430 1370
rect 6464 1368 6520 1370
rect 6554 1368 6631 1370
rect 5669 1349 6631 1368
rect 5669 1345 5741 1349
rect 5669 1311 5688 1345
rect 5722 1311 5741 1345
rect 5669 1255 5741 1311
rect 6559 1326 6631 1349
rect 6559 1292 6578 1326
rect 6612 1292 6631 1326
rect 5669 1221 5688 1255
rect 5722 1221 5741 1255
rect 5669 1165 5741 1221
rect 5669 1131 5688 1165
rect 5722 1131 5741 1165
rect 5669 1075 5741 1131
rect 5669 1041 5688 1075
rect 5722 1041 5741 1075
rect 5669 985 5741 1041
rect 5669 951 5688 985
rect 5722 951 5741 985
rect 5669 895 5741 951
rect 5669 861 5688 895
rect 5722 861 5741 895
rect 5669 805 5741 861
rect 5669 771 5688 805
rect 5722 771 5741 805
rect 5669 715 5741 771
rect 5669 681 5688 715
rect 5722 681 5741 715
rect 5669 625 5741 681
rect 5669 591 5688 625
rect 5722 591 5741 625
rect 5803 1228 6497 1287
rect 5803 1194 5864 1228
rect 5898 1200 5954 1228
rect 5988 1200 6044 1228
rect 6078 1200 6134 1228
rect 5910 1194 5954 1200
rect 6010 1194 6044 1200
rect 6110 1194 6134 1200
rect 6168 1200 6224 1228
rect 6168 1194 6176 1200
rect 5803 1166 5876 1194
rect 5910 1166 5976 1194
rect 6010 1166 6076 1194
rect 6110 1166 6176 1194
rect 6210 1194 6224 1200
rect 6258 1200 6314 1228
rect 6258 1194 6276 1200
rect 6210 1166 6276 1194
rect 6310 1194 6314 1200
rect 6348 1200 6404 1228
rect 6348 1194 6376 1200
rect 6438 1194 6497 1228
rect 6310 1166 6376 1194
rect 6410 1166 6497 1194
rect 5803 1138 6497 1166
rect 5803 1104 5864 1138
rect 5898 1104 5954 1138
rect 5988 1104 6044 1138
rect 6078 1104 6134 1138
rect 6168 1104 6224 1138
rect 6258 1104 6314 1138
rect 6348 1104 6404 1138
rect 6438 1104 6497 1138
rect 5803 1100 6497 1104
rect 5803 1066 5876 1100
rect 5910 1066 5976 1100
rect 6010 1066 6076 1100
rect 6110 1066 6176 1100
rect 6210 1066 6276 1100
rect 6310 1066 6376 1100
rect 6410 1066 6497 1100
rect 5803 1048 6497 1066
rect 5803 1014 5864 1048
rect 5898 1014 5954 1048
rect 5988 1014 6044 1048
rect 6078 1014 6134 1048
rect 6168 1014 6224 1048
rect 6258 1014 6314 1048
rect 6348 1014 6404 1048
rect 6438 1014 6497 1048
rect 5803 1000 6497 1014
rect 5803 966 5876 1000
rect 5910 966 5976 1000
rect 6010 966 6076 1000
rect 6110 966 6176 1000
rect 6210 966 6276 1000
rect 6310 966 6376 1000
rect 6410 966 6497 1000
rect 5803 958 6497 966
rect 5803 924 5864 958
rect 5898 924 5954 958
rect 5988 924 6044 958
rect 6078 924 6134 958
rect 6168 924 6224 958
rect 6258 924 6314 958
rect 6348 924 6404 958
rect 6438 924 6497 958
rect 5803 900 6497 924
rect 5803 868 5876 900
rect 5910 868 5976 900
rect 6010 868 6076 900
rect 6110 868 6176 900
rect 5803 834 5864 868
rect 5910 866 5954 868
rect 6010 866 6044 868
rect 6110 866 6134 868
rect 5898 834 5954 866
rect 5988 834 6044 866
rect 6078 834 6134 866
rect 6168 866 6176 868
rect 6210 868 6276 900
rect 6210 866 6224 868
rect 6168 834 6224 866
rect 6258 866 6276 868
rect 6310 868 6376 900
rect 6410 868 6497 900
rect 6310 866 6314 868
rect 6258 834 6314 866
rect 6348 866 6376 868
rect 6348 834 6404 866
rect 6438 834 6497 868
rect 5803 800 6497 834
rect 5803 778 5876 800
rect 5910 778 5976 800
rect 6010 778 6076 800
rect 6110 778 6176 800
rect 5803 744 5864 778
rect 5910 766 5954 778
rect 6010 766 6044 778
rect 6110 766 6134 778
rect 5898 744 5954 766
rect 5988 744 6044 766
rect 6078 744 6134 766
rect 6168 766 6176 778
rect 6210 778 6276 800
rect 6210 766 6224 778
rect 6168 744 6224 766
rect 6258 766 6276 778
rect 6310 778 6376 800
rect 6410 778 6497 800
rect 6310 766 6314 778
rect 6258 744 6314 766
rect 6348 766 6376 778
rect 6348 744 6404 766
rect 6438 744 6497 778
rect 5803 700 6497 744
rect 5803 688 5876 700
rect 5910 688 5976 700
rect 6010 688 6076 700
rect 6110 688 6176 700
rect 5803 654 5864 688
rect 5910 666 5954 688
rect 6010 666 6044 688
rect 6110 666 6134 688
rect 5898 654 5954 666
rect 5988 654 6044 666
rect 6078 654 6134 666
rect 6168 666 6176 688
rect 6210 688 6276 700
rect 6210 666 6224 688
rect 6168 654 6224 666
rect 6258 666 6276 688
rect 6310 688 6376 700
rect 6410 688 6497 700
rect 6310 666 6314 688
rect 6258 654 6314 666
rect 6348 666 6376 688
rect 6348 654 6404 666
rect 6438 654 6497 688
rect 5803 593 6497 654
rect 6559 1236 6631 1292
rect 6559 1202 6578 1236
rect 6612 1202 6631 1236
rect 6559 1146 6631 1202
rect 6559 1112 6578 1146
rect 6612 1112 6631 1146
rect 6559 1056 6631 1112
rect 6559 1022 6578 1056
rect 6612 1022 6631 1056
rect 6559 966 6631 1022
rect 6559 932 6578 966
rect 6612 932 6631 966
rect 6559 876 6631 932
rect 6559 842 6578 876
rect 6612 842 6631 876
rect 6559 786 6631 842
rect 6559 752 6578 786
rect 6612 752 6631 786
rect 6559 696 6631 752
rect 6559 662 6578 696
rect 6612 662 6631 696
rect 6559 606 6631 662
rect 5669 531 5741 591
rect 6559 572 6578 606
rect 6612 572 6631 606
rect 6559 531 6631 572
rect 5669 512 6631 531
rect 5669 478 5766 512
rect 5800 478 5856 512
rect 5890 478 5946 512
rect 5980 478 6036 512
rect 6070 478 6126 512
rect 6160 478 6216 512
rect 6250 478 6306 512
rect 6340 478 6396 512
rect 6430 478 6486 512
rect 6520 478 6631 512
rect 5669 459 6631 478
rect 6695 1402 6727 1436
rect 6761 1402 6880 1436
rect 6914 1402 6945 1436
rect 8035 1436 8285 1485
rect 6695 1346 6945 1402
rect 6695 1312 6727 1346
rect 6761 1312 6880 1346
rect 6914 1312 6945 1346
rect 6695 1256 6945 1312
rect 6695 1222 6727 1256
rect 6761 1222 6880 1256
rect 6914 1222 6945 1256
rect 6695 1166 6945 1222
rect 6695 1132 6727 1166
rect 6761 1132 6880 1166
rect 6914 1132 6945 1166
rect 6695 1076 6945 1132
rect 6695 1042 6727 1076
rect 6761 1042 6880 1076
rect 6914 1042 6945 1076
rect 6695 986 6945 1042
rect 6695 952 6727 986
rect 6761 952 6880 986
rect 6914 952 6945 986
rect 6695 896 6945 952
rect 6695 862 6727 896
rect 6761 862 6880 896
rect 6914 862 6945 896
rect 6695 806 6945 862
rect 6695 772 6727 806
rect 6761 772 6880 806
rect 6914 772 6945 806
rect 6695 716 6945 772
rect 6695 682 6727 716
rect 6761 682 6880 716
rect 6914 682 6945 716
rect 6695 626 6945 682
rect 6695 592 6727 626
rect 6761 592 6880 626
rect 6914 592 6945 626
rect 6695 536 6945 592
rect 6695 502 6727 536
rect 6761 502 6880 536
rect 6914 502 6945 536
rect 5355 412 5387 446
rect 5421 412 5540 446
rect 5574 412 5605 446
rect 5355 395 5605 412
rect 6695 446 6945 502
rect 7009 1404 7971 1421
rect 7009 1370 7030 1404
rect 7064 1370 7120 1404
rect 7154 1402 7210 1404
rect 7244 1402 7300 1404
rect 7334 1402 7390 1404
rect 7424 1402 7480 1404
rect 7514 1402 7570 1404
rect 7604 1402 7660 1404
rect 7694 1402 7750 1404
rect 7784 1402 7840 1404
rect 7874 1402 7930 1404
rect 7174 1370 7210 1402
rect 7264 1370 7300 1402
rect 7354 1370 7390 1402
rect 7444 1370 7480 1402
rect 7534 1370 7570 1402
rect 7624 1370 7660 1402
rect 7714 1370 7750 1402
rect 7804 1370 7840 1402
rect 7894 1370 7930 1402
rect 7964 1370 7971 1404
rect 7009 1368 7140 1370
rect 7174 1368 7230 1370
rect 7264 1368 7320 1370
rect 7354 1368 7410 1370
rect 7444 1368 7500 1370
rect 7534 1368 7590 1370
rect 7624 1368 7680 1370
rect 7714 1368 7770 1370
rect 7804 1368 7860 1370
rect 7894 1368 7971 1370
rect 7009 1349 7971 1368
rect 7009 1345 7081 1349
rect 7009 1311 7028 1345
rect 7062 1311 7081 1345
rect 7009 1255 7081 1311
rect 7899 1326 7971 1349
rect 7899 1292 7918 1326
rect 7952 1292 7971 1326
rect 7009 1221 7028 1255
rect 7062 1221 7081 1255
rect 7009 1165 7081 1221
rect 7009 1131 7028 1165
rect 7062 1131 7081 1165
rect 7009 1075 7081 1131
rect 7009 1041 7028 1075
rect 7062 1041 7081 1075
rect 7009 985 7081 1041
rect 7009 951 7028 985
rect 7062 951 7081 985
rect 7009 895 7081 951
rect 7009 861 7028 895
rect 7062 861 7081 895
rect 7009 805 7081 861
rect 7009 771 7028 805
rect 7062 771 7081 805
rect 7009 715 7081 771
rect 7009 681 7028 715
rect 7062 681 7081 715
rect 7009 625 7081 681
rect 7009 591 7028 625
rect 7062 591 7081 625
rect 7143 1228 7837 1287
rect 7143 1194 7204 1228
rect 7238 1200 7294 1228
rect 7328 1200 7384 1228
rect 7418 1200 7474 1228
rect 7250 1194 7294 1200
rect 7350 1194 7384 1200
rect 7450 1194 7474 1200
rect 7508 1200 7564 1228
rect 7508 1194 7516 1200
rect 7143 1166 7216 1194
rect 7250 1166 7316 1194
rect 7350 1166 7416 1194
rect 7450 1166 7516 1194
rect 7550 1194 7564 1200
rect 7598 1200 7654 1228
rect 7598 1194 7616 1200
rect 7550 1166 7616 1194
rect 7650 1194 7654 1200
rect 7688 1200 7744 1228
rect 7688 1194 7716 1200
rect 7778 1194 7837 1228
rect 7650 1166 7716 1194
rect 7750 1166 7837 1194
rect 7143 1138 7837 1166
rect 7143 1104 7204 1138
rect 7238 1104 7294 1138
rect 7328 1104 7384 1138
rect 7418 1104 7474 1138
rect 7508 1104 7564 1138
rect 7598 1104 7654 1138
rect 7688 1104 7744 1138
rect 7778 1104 7837 1138
rect 7143 1100 7837 1104
rect 7143 1066 7216 1100
rect 7250 1066 7316 1100
rect 7350 1066 7416 1100
rect 7450 1066 7516 1100
rect 7550 1066 7616 1100
rect 7650 1066 7716 1100
rect 7750 1066 7837 1100
rect 7143 1048 7837 1066
rect 7143 1014 7204 1048
rect 7238 1014 7294 1048
rect 7328 1014 7384 1048
rect 7418 1014 7474 1048
rect 7508 1014 7564 1048
rect 7598 1014 7654 1048
rect 7688 1014 7744 1048
rect 7778 1014 7837 1048
rect 7143 1000 7837 1014
rect 7143 966 7216 1000
rect 7250 966 7316 1000
rect 7350 966 7416 1000
rect 7450 966 7516 1000
rect 7550 966 7616 1000
rect 7650 966 7716 1000
rect 7750 966 7837 1000
rect 7143 958 7837 966
rect 7143 924 7204 958
rect 7238 924 7294 958
rect 7328 924 7384 958
rect 7418 924 7474 958
rect 7508 924 7564 958
rect 7598 924 7654 958
rect 7688 924 7744 958
rect 7778 924 7837 958
rect 7143 900 7837 924
rect 7143 868 7216 900
rect 7250 868 7316 900
rect 7350 868 7416 900
rect 7450 868 7516 900
rect 7143 834 7204 868
rect 7250 866 7294 868
rect 7350 866 7384 868
rect 7450 866 7474 868
rect 7238 834 7294 866
rect 7328 834 7384 866
rect 7418 834 7474 866
rect 7508 866 7516 868
rect 7550 868 7616 900
rect 7550 866 7564 868
rect 7508 834 7564 866
rect 7598 866 7616 868
rect 7650 868 7716 900
rect 7750 868 7837 900
rect 7650 866 7654 868
rect 7598 834 7654 866
rect 7688 866 7716 868
rect 7688 834 7744 866
rect 7778 834 7837 868
rect 7143 800 7837 834
rect 7143 778 7216 800
rect 7250 778 7316 800
rect 7350 778 7416 800
rect 7450 778 7516 800
rect 7143 744 7204 778
rect 7250 766 7294 778
rect 7350 766 7384 778
rect 7450 766 7474 778
rect 7238 744 7294 766
rect 7328 744 7384 766
rect 7418 744 7474 766
rect 7508 766 7516 778
rect 7550 778 7616 800
rect 7550 766 7564 778
rect 7508 744 7564 766
rect 7598 766 7616 778
rect 7650 778 7716 800
rect 7750 778 7837 800
rect 7650 766 7654 778
rect 7598 744 7654 766
rect 7688 766 7716 778
rect 7688 744 7744 766
rect 7778 744 7837 778
rect 7143 700 7837 744
rect 7143 688 7216 700
rect 7250 688 7316 700
rect 7350 688 7416 700
rect 7450 688 7516 700
rect 7143 654 7204 688
rect 7250 666 7294 688
rect 7350 666 7384 688
rect 7450 666 7474 688
rect 7238 654 7294 666
rect 7328 654 7384 666
rect 7418 654 7474 666
rect 7508 666 7516 688
rect 7550 688 7616 700
rect 7550 666 7564 688
rect 7508 654 7564 666
rect 7598 666 7616 688
rect 7650 688 7716 700
rect 7750 688 7837 700
rect 7650 666 7654 688
rect 7598 654 7654 666
rect 7688 666 7716 688
rect 7688 654 7744 666
rect 7778 654 7837 688
rect 7143 593 7837 654
rect 7899 1236 7971 1292
rect 7899 1202 7918 1236
rect 7952 1202 7971 1236
rect 7899 1146 7971 1202
rect 7899 1112 7918 1146
rect 7952 1112 7971 1146
rect 7899 1056 7971 1112
rect 7899 1022 7918 1056
rect 7952 1022 7971 1056
rect 7899 966 7971 1022
rect 7899 932 7918 966
rect 7952 932 7971 966
rect 7899 876 7971 932
rect 7899 842 7918 876
rect 7952 842 7971 876
rect 7899 786 7971 842
rect 7899 752 7918 786
rect 7952 752 7971 786
rect 7899 696 7971 752
rect 7899 662 7918 696
rect 7952 662 7971 696
rect 7899 606 7971 662
rect 7009 531 7081 591
rect 7899 572 7918 606
rect 7952 572 7971 606
rect 7899 531 7971 572
rect 7009 512 7971 531
rect 7009 478 7106 512
rect 7140 478 7196 512
rect 7230 478 7286 512
rect 7320 478 7376 512
rect 7410 478 7466 512
rect 7500 478 7556 512
rect 7590 478 7646 512
rect 7680 478 7736 512
rect 7770 478 7826 512
rect 7860 478 7971 512
rect 7009 459 7971 478
rect 8035 1402 8067 1436
rect 8101 1402 8220 1436
rect 8254 1402 8285 1436
rect 9375 1436 9625 1485
rect 8035 1346 8285 1402
rect 8035 1312 8067 1346
rect 8101 1312 8220 1346
rect 8254 1312 8285 1346
rect 8035 1256 8285 1312
rect 8035 1222 8067 1256
rect 8101 1222 8220 1256
rect 8254 1222 8285 1256
rect 8035 1166 8285 1222
rect 8035 1132 8067 1166
rect 8101 1132 8220 1166
rect 8254 1132 8285 1166
rect 8035 1076 8285 1132
rect 8035 1042 8067 1076
rect 8101 1042 8220 1076
rect 8254 1042 8285 1076
rect 8035 986 8285 1042
rect 8035 952 8067 986
rect 8101 952 8220 986
rect 8254 952 8285 986
rect 8035 896 8285 952
rect 8035 862 8067 896
rect 8101 862 8220 896
rect 8254 862 8285 896
rect 8035 806 8285 862
rect 8035 772 8067 806
rect 8101 772 8220 806
rect 8254 772 8285 806
rect 8035 716 8285 772
rect 8035 682 8067 716
rect 8101 682 8220 716
rect 8254 682 8285 716
rect 8035 626 8285 682
rect 8035 592 8067 626
rect 8101 592 8220 626
rect 8254 592 8285 626
rect 8035 536 8285 592
rect 8035 502 8067 536
rect 8101 502 8220 536
rect 8254 502 8285 536
rect 6695 412 6727 446
rect 6761 412 6880 446
rect 6914 412 6945 446
rect 6695 395 6945 412
rect 8035 446 8285 502
rect 8349 1404 9311 1421
rect 8349 1370 8370 1404
rect 8404 1370 8460 1404
rect 8494 1402 8550 1404
rect 8584 1402 8640 1404
rect 8674 1402 8730 1404
rect 8764 1402 8820 1404
rect 8854 1402 8910 1404
rect 8944 1402 9000 1404
rect 9034 1402 9090 1404
rect 9124 1402 9180 1404
rect 9214 1402 9270 1404
rect 8514 1370 8550 1402
rect 8604 1370 8640 1402
rect 8694 1370 8730 1402
rect 8784 1370 8820 1402
rect 8874 1370 8910 1402
rect 8964 1370 9000 1402
rect 9054 1370 9090 1402
rect 9144 1370 9180 1402
rect 9234 1370 9270 1402
rect 9304 1370 9311 1404
rect 8349 1368 8480 1370
rect 8514 1368 8570 1370
rect 8604 1368 8660 1370
rect 8694 1368 8750 1370
rect 8784 1368 8840 1370
rect 8874 1368 8930 1370
rect 8964 1368 9020 1370
rect 9054 1368 9110 1370
rect 9144 1368 9200 1370
rect 9234 1368 9311 1370
rect 8349 1349 9311 1368
rect 8349 1345 8421 1349
rect 8349 1311 8368 1345
rect 8402 1311 8421 1345
rect 8349 1255 8421 1311
rect 9239 1326 9311 1349
rect 9239 1292 9258 1326
rect 9292 1292 9311 1326
rect 8349 1221 8368 1255
rect 8402 1221 8421 1255
rect 8349 1165 8421 1221
rect 8349 1131 8368 1165
rect 8402 1131 8421 1165
rect 8349 1075 8421 1131
rect 8349 1041 8368 1075
rect 8402 1041 8421 1075
rect 8349 985 8421 1041
rect 8349 951 8368 985
rect 8402 951 8421 985
rect 8349 895 8421 951
rect 8349 861 8368 895
rect 8402 861 8421 895
rect 8349 805 8421 861
rect 8349 771 8368 805
rect 8402 771 8421 805
rect 8349 715 8421 771
rect 8349 681 8368 715
rect 8402 681 8421 715
rect 8349 625 8421 681
rect 8349 591 8368 625
rect 8402 591 8421 625
rect 8483 1228 9177 1287
rect 8483 1194 8544 1228
rect 8578 1200 8634 1228
rect 8668 1200 8724 1228
rect 8758 1200 8814 1228
rect 8590 1194 8634 1200
rect 8690 1194 8724 1200
rect 8790 1194 8814 1200
rect 8848 1200 8904 1228
rect 8848 1194 8856 1200
rect 8483 1166 8556 1194
rect 8590 1166 8656 1194
rect 8690 1166 8756 1194
rect 8790 1166 8856 1194
rect 8890 1194 8904 1200
rect 8938 1200 8994 1228
rect 8938 1194 8956 1200
rect 8890 1166 8956 1194
rect 8990 1194 8994 1200
rect 9028 1200 9084 1228
rect 9028 1194 9056 1200
rect 9118 1194 9177 1228
rect 8990 1166 9056 1194
rect 9090 1166 9177 1194
rect 8483 1138 9177 1166
rect 8483 1104 8544 1138
rect 8578 1104 8634 1138
rect 8668 1104 8724 1138
rect 8758 1104 8814 1138
rect 8848 1104 8904 1138
rect 8938 1104 8994 1138
rect 9028 1104 9084 1138
rect 9118 1104 9177 1138
rect 8483 1100 9177 1104
rect 8483 1066 8556 1100
rect 8590 1066 8656 1100
rect 8690 1066 8756 1100
rect 8790 1066 8856 1100
rect 8890 1066 8956 1100
rect 8990 1066 9056 1100
rect 9090 1066 9177 1100
rect 8483 1048 9177 1066
rect 8483 1014 8544 1048
rect 8578 1014 8634 1048
rect 8668 1014 8724 1048
rect 8758 1014 8814 1048
rect 8848 1014 8904 1048
rect 8938 1014 8994 1048
rect 9028 1014 9084 1048
rect 9118 1014 9177 1048
rect 8483 1000 9177 1014
rect 8483 966 8556 1000
rect 8590 966 8656 1000
rect 8690 966 8756 1000
rect 8790 966 8856 1000
rect 8890 966 8956 1000
rect 8990 966 9056 1000
rect 9090 966 9177 1000
rect 8483 958 9177 966
rect 8483 924 8544 958
rect 8578 924 8634 958
rect 8668 924 8724 958
rect 8758 924 8814 958
rect 8848 924 8904 958
rect 8938 924 8994 958
rect 9028 924 9084 958
rect 9118 924 9177 958
rect 8483 900 9177 924
rect 8483 868 8556 900
rect 8590 868 8656 900
rect 8690 868 8756 900
rect 8790 868 8856 900
rect 8483 834 8544 868
rect 8590 866 8634 868
rect 8690 866 8724 868
rect 8790 866 8814 868
rect 8578 834 8634 866
rect 8668 834 8724 866
rect 8758 834 8814 866
rect 8848 866 8856 868
rect 8890 868 8956 900
rect 8890 866 8904 868
rect 8848 834 8904 866
rect 8938 866 8956 868
rect 8990 868 9056 900
rect 9090 868 9177 900
rect 8990 866 8994 868
rect 8938 834 8994 866
rect 9028 866 9056 868
rect 9028 834 9084 866
rect 9118 834 9177 868
rect 8483 800 9177 834
rect 8483 778 8556 800
rect 8590 778 8656 800
rect 8690 778 8756 800
rect 8790 778 8856 800
rect 8483 744 8544 778
rect 8590 766 8634 778
rect 8690 766 8724 778
rect 8790 766 8814 778
rect 8578 744 8634 766
rect 8668 744 8724 766
rect 8758 744 8814 766
rect 8848 766 8856 778
rect 8890 778 8956 800
rect 8890 766 8904 778
rect 8848 744 8904 766
rect 8938 766 8956 778
rect 8990 778 9056 800
rect 9090 778 9177 800
rect 8990 766 8994 778
rect 8938 744 8994 766
rect 9028 766 9056 778
rect 9028 744 9084 766
rect 9118 744 9177 778
rect 8483 700 9177 744
rect 8483 688 8556 700
rect 8590 688 8656 700
rect 8690 688 8756 700
rect 8790 688 8856 700
rect 8483 654 8544 688
rect 8590 666 8634 688
rect 8690 666 8724 688
rect 8790 666 8814 688
rect 8578 654 8634 666
rect 8668 654 8724 666
rect 8758 654 8814 666
rect 8848 666 8856 688
rect 8890 688 8956 700
rect 8890 666 8904 688
rect 8848 654 8904 666
rect 8938 666 8956 688
rect 8990 688 9056 700
rect 9090 688 9177 700
rect 8990 666 8994 688
rect 8938 654 8994 666
rect 9028 666 9056 688
rect 9028 654 9084 666
rect 9118 654 9177 688
rect 8483 593 9177 654
rect 9239 1236 9311 1292
rect 9239 1202 9258 1236
rect 9292 1202 9311 1236
rect 9239 1146 9311 1202
rect 9239 1112 9258 1146
rect 9292 1112 9311 1146
rect 9239 1056 9311 1112
rect 9239 1022 9258 1056
rect 9292 1022 9311 1056
rect 9239 966 9311 1022
rect 9239 932 9258 966
rect 9292 932 9311 966
rect 9239 876 9311 932
rect 9239 842 9258 876
rect 9292 842 9311 876
rect 9239 786 9311 842
rect 9239 752 9258 786
rect 9292 752 9311 786
rect 9239 696 9311 752
rect 9239 662 9258 696
rect 9292 662 9311 696
rect 9239 606 9311 662
rect 8349 531 8421 591
rect 9239 572 9258 606
rect 9292 572 9311 606
rect 9239 531 9311 572
rect 8349 512 9311 531
rect 8349 478 8446 512
rect 8480 478 8536 512
rect 8570 478 8626 512
rect 8660 478 8716 512
rect 8750 478 8806 512
rect 8840 478 8896 512
rect 8930 478 8986 512
rect 9020 478 9076 512
rect 9110 478 9166 512
rect 9200 478 9311 512
rect 8349 459 9311 478
rect 9375 1402 9407 1436
rect 9441 1402 9560 1436
rect 9594 1402 9625 1436
rect 10715 1436 10814 1485
rect 9375 1346 9625 1402
rect 9375 1312 9407 1346
rect 9441 1312 9560 1346
rect 9594 1312 9625 1346
rect 9375 1256 9625 1312
rect 9375 1222 9407 1256
rect 9441 1222 9560 1256
rect 9594 1222 9625 1256
rect 9375 1166 9625 1222
rect 9375 1132 9407 1166
rect 9441 1132 9560 1166
rect 9594 1132 9625 1166
rect 9375 1076 9625 1132
rect 9375 1042 9407 1076
rect 9441 1042 9560 1076
rect 9594 1042 9625 1076
rect 9375 986 9625 1042
rect 9375 952 9407 986
rect 9441 952 9560 986
rect 9594 952 9625 986
rect 9375 896 9625 952
rect 9375 862 9407 896
rect 9441 862 9560 896
rect 9594 862 9625 896
rect 9375 806 9625 862
rect 9375 772 9407 806
rect 9441 772 9560 806
rect 9594 772 9625 806
rect 9375 716 9625 772
rect 9375 682 9407 716
rect 9441 682 9560 716
rect 9594 682 9625 716
rect 9375 626 9625 682
rect 9375 592 9407 626
rect 9441 592 9560 626
rect 9594 592 9625 626
rect 9375 536 9625 592
rect 9375 502 9407 536
rect 9441 502 9560 536
rect 9594 502 9625 536
rect 8035 412 8067 446
rect 8101 412 8220 446
rect 8254 412 8285 446
rect 8035 395 8285 412
rect 9375 446 9625 502
rect 9689 1404 10651 1421
rect 9689 1370 9710 1404
rect 9744 1370 9800 1404
rect 9834 1402 9890 1404
rect 9924 1402 9980 1404
rect 10014 1402 10070 1404
rect 10104 1402 10160 1404
rect 10194 1402 10250 1404
rect 10284 1402 10340 1404
rect 10374 1402 10430 1404
rect 10464 1402 10520 1404
rect 10554 1402 10610 1404
rect 9854 1370 9890 1402
rect 9944 1370 9980 1402
rect 10034 1370 10070 1402
rect 10124 1370 10160 1402
rect 10214 1370 10250 1402
rect 10304 1370 10340 1402
rect 10394 1370 10430 1402
rect 10484 1370 10520 1402
rect 10574 1370 10610 1402
rect 10644 1370 10651 1404
rect 9689 1368 9820 1370
rect 9854 1368 9910 1370
rect 9944 1368 10000 1370
rect 10034 1368 10090 1370
rect 10124 1368 10180 1370
rect 10214 1368 10270 1370
rect 10304 1368 10360 1370
rect 10394 1368 10450 1370
rect 10484 1368 10540 1370
rect 10574 1368 10651 1370
rect 9689 1349 10651 1368
rect 9689 1345 9761 1349
rect 9689 1311 9708 1345
rect 9742 1311 9761 1345
rect 9689 1255 9761 1311
rect 10579 1326 10651 1349
rect 10579 1292 10598 1326
rect 10632 1292 10651 1326
rect 9689 1221 9708 1255
rect 9742 1221 9761 1255
rect 9689 1165 9761 1221
rect 9689 1131 9708 1165
rect 9742 1131 9761 1165
rect 9689 1075 9761 1131
rect 9689 1041 9708 1075
rect 9742 1041 9761 1075
rect 9689 985 9761 1041
rect 9689 951 9708 985
rect 9742 951 9761 985
rect 9689 895 9761 951
rect 9689 861 9708 895
rect 9742 861 9761 895
rect 9689 805 9761 861
rect 9689 771 9708 805
rect 9742 771 9761 805
rect 9689 715 9761 771
rect 9689 681 9708 715
rect 9742 681 9761 715
rect 9689 625 9761 681
rect 9689 591 9708 625
rect 9742 591 9761 625
rect 9823 1228 10517 1287
rect 9823 1194 9884 1228
rect 9918 1200 9974 1228
rect 10008 1200 10064 1228
rect 10098 1200 10154 1228
rect 9930 1194 9974 1200
rect 10030 1194 10064 1200
rect 10130 1194 10154 1200
rect 10188 1200 10244 1228
rect 10188 1194 10196 1200
rect 9823 1166 9896 1194
rect 9930 1166 9996 1194
rect 10030 1166 10096 1194
rect 10130 1166 10196 1194
rect 10230 1194 10244 1200
rect 10278 1200 10334 1228
rect 10278 1194 10296 1200
rect 10230 1166 10296 1194
rect 10330 1194 10334 1200
rect 10368 1200 10424 1228
rect 10368 1194 10396 1200
rect 10458 1194 10517 1228
rect 10330 1166 10396 1194
rect 10430 1166 10517 1194
rect 9823 1138 10517 1166
rect 9823 1104 9884 1138
rect 9918 1104 9974 1138
rect 10008 1104 10064 1138
rect 10098 1104 10154 1138
rect 10188 1104 10244 1138
rect 10278 1104 10334 1138
rect 10368 1104 10424 1138
rect 10458 1104 10517 1138
rect 9823 1100 10517 1104
rect 9823 1066 9896 1100
rect 9930 1066 9996 1100
rect 10030 1066 10096 1100
rect 10130 1066 10196 1100
rect 10230 1066 10296 1100
rect 10330 1066 10396 1100
rect 10430 1066 10517 1100
rect 9823 1048 10517 1066
rect 9823 1014 9884 1048
rect 9918 1014 9974 1048
rect 10008 1014 10064 1048
rect 10098 1014 10154 1048
rect 10188 1014 10244 1048
rect 10278 1014 10334 1048
rect 10368 1014 10424 1048
rect 10458 1014 10517 1048
rect 9823 1000 10517 1014
rect 9823 966 9896 1000
rect 9930 966 9996 1000
rect 10030 966 10096 1000
rect 10130 966 10196 1000
rect 10230 966 10296 1000
rect 10330 966 10396 1000
rect 10430 966 10517 1000
rect 9823 958 10517 966
rect 9823 924 9884 958
rect 9918 924 9974 958
rect 10008 924 10064 958
rect 10098 924 10154 958
rect 10188 924 10244 958
rect 10278 924 10334 958
rect 10368 924 10424 958
rect 10458 924 10517 958
rect 9823 900 10517 924
rect 9823 868 9896 900
rect 9930 868 9996 900
rect 10030 868 10096 900
rect 10130 868 10196 900
rect 9823 834 9884 868
rect 9930 866 9974 868
rect 10030 866 10064 868
rect 10130 866 10154 868
rect 9918 834 9974 866
rect 10008 834 10064 866
rect 10098 834 10154 866
rect 10188 866 10196 868
rect 10230 868 10296 900
rect 10230 866 10244 868
rect 10188 834 10244 866
rect 10278 866 10296 868
rect 10330 868 10396 900
rect 10430 868 10517 900
rect 10330 866 10334 868
rect 10278 834 10334 866
rect 10368 866 10396 868
rect 10368 834 10424 866
rect 10458 834 10517 868
rect 9823 800 10517 834
rect 9823 778 9896 800
rect 9930 778 9996 800
rect 10030 778 10096 800
rect 10130 778 10196 800
rect 9823 744 9884 778
rect 9930 766 9974 778
rect 10030 766 10064 778
rect 10130 766 10154 778
rect 9918 744 9974 766
rect 10008 744 10064 766
rect 10098 744 10154 766
rect 10188 766 10196 778
rect 10230 778 10296 800
rect 10230 766 10244 778
rect 10188 744 10244 766
rect 10278 766 10296 778
rect 10330 778 10396 800
rect 10430 778 10517 800
rect 10330 766 10334 778
rect 10278 744 10334 766
rect 10368 766 10396 778
rect 10368 744 10424 766
rect 10458 744 10517 778
rect 9823 700 10517 744
rect 9823 688 9896 700
rect 9930 688 9996 700
rect 10030 688 10096 700
rect 10130 688 10196 700
rect 9823 654 9884 688
rect 9930 666 9974 688
rect 10030 666 10064 688
rect 10130 666 10154 688
rect 9918 654 9974 666
rect 10008 654 10064 666
rect 10098 654 10154 666
rect 10188 666 10196 688
rect 10230 688 10296 700
rect 10230 666 10244 688
rect 10188 654 10244 666
rect 10278 666 10296 688
rect 10330 688 10396 700
rect 10430 688 10517 700
rect 10330 666 10334 688
rect 10278 654 10334 666
rect 10368 666 10396 688
rect 10368 654 10424 666
rect 10458 654 10517 688
rect 9823 593 10517 654
rect 10579 1236 10651 1292
rect 10579 1202 10598 1236
rect 10632 1202 10651 1236
rect 10579 1146 10651 1202
rect 10579 1112 10598 1146
rect 10632 1112 10651 1146
rect 10579 1056 10651 1112
rect 10579 1022 10598 1056
rect 10632 1022 10651 1056
rect 10579 966 10651 1022
rect 10579 932 10598 966
rect 10632 932 10651 966
rect 10579 876 10651 932
rect 10579 842 10598 876
rect 10632 842 10651 876
rect 10579 786 10651 842
rect 10579 752 10598 786
rect 10632 752 10651 786
rect 10579 696 10651 752
rect 10579 662 10598 696
rect 10632 662 10651 696
rect 10579 606 10651 662
rect 9689 531 9761 591
rect 10579 572 10598 606
rect 10632 572 10651 606
rect 10579 531 10651 572
rect 9689 512 10651 531
rect 9689 478 9786 512
rect 9820 478 9876 512
rect 9910 478 9966 512
rect 10000 478 10056 512
rect 10090 478 10146 512
rect 10180 478 10236 512
rect 10270 478 10326 512
rect 10360 478 10416 512
rect 10450 478 10506 512
rect 10540 478 10651 512
rect 9689 459 10651 478
rect 10715 1402 10747 1436
rect 10781 1402 10814 1436
rect 10715 1346 10814 1402
rect 10715 1312 10747 1346
rect 10781 1312 10814 1346
rect 10715 1256 10814 1312
rect 10715 1222 10747 1256
rect 10781 1222 10814 1256
rect 10715 1166 10814 1222
rect 10715 1132 10747 1166
rect 10781 1132 10814 1166
rect 10715 1076 10814 1132
rect 10715 1042 10747 1076
rect 10781 1042 10814 1076
rect 10715 986 10814 1042
rect 10715 952 10747 986
rect 10781 952 10814 986
rect 10715 896 10814 952
rect 10715 862 10747 896
rect 10781 862 10814 896
rect 10715 806 10814 862
rect 10715 772 10747 806
rect 10781 772 10814 806
rect 10715 716 10814 772
rect 10715 682 10747 716
rect 10781 682 10814 716
rect 10715 626 10814 682
rect 10715 592 10747 626
rect 10781 592 10814 626
rect 10715 536 10814 592
rect 10715 502 10747 536
rect 10781 502 10814 536
rect 9375 412 9407 446
rect 9441 412 9560 446
rect 9594 412 9625 446
rect 9375 395 9625 412
rect 10715 446 10814 502
rect 10715 412 10747 446
rect 10781 412 10814 446
rect 10715 395 10814 412
rect 146 362 10814 395
rect 146 328 276 362
rect 310 328 366 362
rect 400 328 456 362
rect 490 328 546 362
rect 580 328 636 362
rect 670 328 726 362
rect 760 328 816 362
rect 850 328 906 362
rect 940 328 996 362
rect 1030 328 1086 362
rect 1120 328 1176 362
rect 1210 328 1266 362
rect 1300 328 1616 362
rect 1650 328 1706 362
rect 1740 328 1796 362
rect 1830 328 1886 362
rect 1920 328 1976 362
rect 2010 328 2066 362
rect 2100 328 2156 362
rect 2190 328 2246 362
rect 2280 328 2336 362
rect 2370 328 2426 362
rect 2460 328 2516 362
rect 2550 328 2606 362
rect 2640 328 2956 362
rect 2990 328 3046 362
rect 3080 328 3136 362
rect 3170 328 3226 362
rect 3260 328 3316 362
rect 3350 328 3406 362
rect 3440 328 3496 362
rect 3530 328 3586 362
rect 3620 328 3676 362
rect 3710 328 3766 362
rect 3800 328 3856 362
rect 3890 328 3946 362
rect 3980 328 4296 362
rect 4330 328 4386 362
rect 4420 328 4476 362
rect 4510 328 4566 362
rect 4600 328 4656 362
rect 4690 328 4746 362
rect 4780 328 4836 362
rect 4870 328 4926 362
rect 4960 328 5016 362
rect 5050 328 5106 362
rect 5140 328 5196 362
rect 5230 328 5286 362
rect 5320 328 5636 362
rect 5670 328 5726 362
rect 5760 328 5816 362
rect 5850 328 5906 362
rect 5940 328 5996 362
rect 6030 328 6086 362
rect 6120 328 6176 362
rect 6210 328 6266 362
rect 6300 328 6356 362
rect 6390 328 6446 362
rect 6480 328 6536 362
rect 6570 328 6626 362
rect 6660 328 6976 362
rect 7010 328 7066 362
rect 7100 328 7156 362
rect 7190 328 7246 362
rect 7280 328 7336 362
rect 7370 328 7426 362
rect 7460 328 7516 362
rect 7550 328 7606 362
rect 7640 328 7696 362
rect 7730 328 7786 362
rect 7820 328 7876 362
rect 7910 328 7966 362
rect 8000 328 8316 362
rect 8350 328 8406 362
rect 8440 328 8496 362
rect 8530 328 8586 362
rect 8620 328 8676 362
rect 8710 328 8766 362
rect 8800 328 8856 362
rect 8890 328 8946 362
rect 8980 328 9036 362
rect 9070 328 9126 362
rect 9160 328 9216 362
rect 9250 328 9306 362
rect 9340 328 9656 362
rect 9690 328 9746 362
rect 9780 328 9836 362
rect 9870 328 9926 362
rect 9960 328 10016 362
rect 10050 328 10106 362
rect 10140 328 10196 362
rect 10230 328 10286 362
rect 10320 328 10376 362
rect 10410 328 10466 362
rect 10500 328 10556 362
rect 10590 328 10646 362
rect 10680 328 10814 362
rect 146 296 10814 328
rect 120 17 10840 30
rect 120 -17 303 17
rect 337 -17 503 17
rect 537 -17 703 17
rect 737 -17 903 17
rect 937 -17 1103 17
rect 1137 -17 1303 17
rect 1337 -17 1503 17
rect 1537 -17 1703 17
rect 1737 -17 1903 17
rect 1937 -17 2103 17
rect 2137 -17 2303 17
rect 2337 -17 2503 17
rect 2537 -17 2703 17
rect 2737 -17 2903 17
rect 2937 -17 3103 17
rect 3137 -17 3303 17
rect 3337 -17 3503 17
rect 3537 -17 3703 17
rect 3737 -17 3903 17
rect 3937 -17 4103 17
rect 4137 -17 4303 17
rect 4337 -17 4503 17
rect 4537 -17 4703 17
rect 4737 -17 4903 17
rect 4937 -17 5103 17
rect 5137 -17 5303 17
rect 5337 -17 5503 17
rect 5537 -17 5703 17
rect 5737 -17 5903 17
rect 5937 -17 6103 17
rect 6137 -17 6303 17
rect 6337 -17 6503 17
rect 6537 -17 6703 17
rect 6737 -17 6903 17
rect 6937 -17 7103 17
rect 7137 -17 7303 17
rect 7337 -17 7503 17
rect 7537 -17 7703 17
rect 7737 -17 7903 17
rect 7937 -17 8103 17
rect 8137 -17 8303 17
rect 8337 -17 8503 17
rect 8537 -17 8703 17
rect 8737 -17 8903 17
rect 8937 -17 9103 17
rect 9137 -17 9303 17
rect 9337 -17 9503 17
rect 9537 -17 9703 17
rect 9737 -17 9903 17
rect 9937 -17 10103 17
rect 10137 -17 10303 17
rect 10337 -17 10503 17
rect 10537 -17 10703 17
rect 10737 -17 10840 17
rect 120 -30 10840 -17
<< viali >>
rect 303 1863 337 1897
rect 503 1863 537 1897
rect 703 1863 737 1897
rect 903 1863 937 1897
rect 1103 1863 1137 1897
rect 1303 1863 1337 1897
rect 1503 1863 1537 1897
rect 1703 1863 1737 1897
rect 1903 1863 1937 1897
rect 2103 1863 2137 1897
rect 2303 1863 2337 1897
rect 2503 1863 2537 1897
rect 2703 1863 2737 1897
rect 2903 1863 2937 1897
rect 3103 1863 3137 1897
rect 3303 1863 3337 1897
rect 3503 1863 3537 1897
rect 3703 1863 3737 1897
rect 3903 1863 3937 1897
rect 4103 1863 4137 1897
rect 4303 1863 4337 1897
rect 4503 1863 4537 1897
rect 4703 1863 4737 1897
rect 4903 1863 4937 1897
rect 5103 1863 5137 1897
rect 5303 1863 5337 1897
rect 5503 1863 5537 1897
rect 5703 1863 5737 1897
rect 5903 1863 5937 1897
rect 6103 1863 6137 1897
rect 6303 1863 6337 1897
rect 6503 1863 6537 1897
rect 6703 1863 6737 1897
rect 6903 1863 6937 1897
rect 7103 1863 7137 1897
rect 7303 1863 7337 1897
rect 7503 1863 7537 1897
rect 7703 1863 7737 1897
rect 7903 1863 7937 1897
rect 8103 1863 8137 1897
rect 8303 1863 8337 1897
rect 8503 1863 8537 1897
rect 8703 1863 8737 1897
rect 8903 1863 8937 1897
rect 9103 1863 9137 1897
rect 9303 1863 9337 1897
rect 9503 1863 9537 1897
rect 9703 1863 9737 1897
rect 9903 1863 9937 1897
rect 10103 1863 10137 1897
rect 10303 1863 10337 1897
rect 10503 1863 10537 1897
rect 10703 1863 10737 1897
rect 166 1530 200 1564
rect 256 1549 290 1564
rect 346 1549 380 1564
rect 436 1549 470 1564
rect 526 1549 560 1564
rect 616 1549 650 1564
rect 706 1549 740 1564
rect 796 1549 830 1564
rect 886 1549 920 1564
rect 976 1549 1010 1564
rect 1066 1549 1100 1564
rect 1156 1549 1190 1564
rect 1246 1549 1280 1564
rect 256 1530 276 1549
rect 276 1530 290 1549
rect 346 1530 366 1549
rect 366 1530 380 1549
rect 436 1530 456 1549
rect 456 1530 470 1549
rect 526 1530 546 1549
rect 546 1530 560 1549
rect 616 1530 636 1549
rect 636 1530 650 1549
rect 706 1530 726 1549
rect 726 1530 740 1549
rect 796 1530 816 1549
rect 816 1530 830 1549
rect 886 1530 906 1549
rect 906 1530 920 1549
rect 976 1530 996 1549
rect 996 1530 1010 1549
rect 1066 1530 1086 1549
rect 1086 1530 1100 1549
rect 1156 1530 1176 1549
rect 1176 1530 1190 1549
rect 1246 1530 1266 1549
rect 1266 1530 1280 1549
rect 1336 1530 1370 1564
rect 1506 1530 1540 1564
rect 1596 1549 1630 1564
rect 1686 1549 1720 1564
rect 1776 1549 1810 1564
rect 1866 1549 1900 1564
rect 1956 1549 1990 1564
rect 2046 1549 2080 1564
rect 2136 1549 2170 1564
rect 2226 1549 2260 1564
rect 2316 1549 2350 1564
rect 2406 1549 2440 1564
rect 2496 1549 2530 1564
rect 2586 1549 2620 1564
rect 1596 1530 1616 1549
rect 1616 1530 1630 1549
rect 1686 1530 1706 1549
rect 1706 1530 1720 1549
rect 1776 1530 1796 1549
rect 1796 1530 1810 1549
rect 1866 1530 1886 1549
rect 1886 1530 1900 1549
rect 1956 1530 1976 1549
rect 1976 1530 1990 1549
rect 2046 1530 2066 1549
rect 2066 1530 2080 1549
rect 2136 1530 2156 1549
rect 2156 1530 2170 1549
rect 2226 1530 2246 1549
rect 2246 1530 2260 1549
rect 2316 1530 2336 1549
rect 2336 1530 2350 1549
rect 2406 1530 2426 1549
rect 2426 1530 2440 1549
rect 2496 1530 2516 1549
rect 2516 1530 2530 1549
rect 2586 1530 2606 1549
rect 2606 1530 2620 1549
rect 2676 1530 2710 1564
rect 2846 1530 2880 1564
rect 2936 1549 2970 1564
rect 3026 1549 3060 1564
rect 3116 1549 3150 1564
rect 3206 1549 3240 1564
rect 3296 1549 3330 1564
rect 3386 1549 3420 1564
rect 3476 1549 3510 1564
rect 3566 1549 3600 1564
rect 3656 1549 3690 1564
rect 3746 1549 3780 1564
rect 3836 1549 3870 1564
rect 3926 1549 3960 1564
rect 2936 1530 2956 1549
rect 2956 1530 2970 1549
rect 3026 1530 3046 1549
rect 3046 1530 3060 1549
rect 3116 1530 3136 1549
rect 3136 1530 3150 1549
rect 3206 1530 3226 1549
rect 3226 1530 3240 1549
rect 3296 1530 3316 1549
rect 3316 1530 3330 1549
rect 3386 1530 3406 1549
rect 3406 1530 3420 1549
rect 3476 1530 3496 1549
rect 3496 1530 3510 1549
rect 3566 1530 3586 1549
rect 3586 1530 3600 1549
rect 3656 1530 3676 1549
rect 3676 1530 3690 1549
rect 3746 1530 3766 1549
rect 3766 1530 3780 1549
rect 3836 1530 3856 1549
rect 3856 1530 3870 1549
rect 3926 1530 3946 1549
rect 3946 1530 3960 1549
rect 4016 1530 4050 1564
rect 4186 1530 4220 1564
rect 4276 1549 4310 1564
rect 4366 1549 4400 1564
rect 4456 1549 4490 1564
rect 4546 1549 4580 1564
rect 4636 1549 4670 1564
rect 4726 1549 4760 1564
rect 4816 1549 4850 1564
rect 4906 1549 4940 1564
rect 4996 1549 5030 1564
rect 5086 1549 5120 1564
rect 5176 1549 5210 1564
rect 5266 1549 5300 1564
rect 4276 1530 4296 1549
rect 4296 1530 4310 1549
rect 4366 1530 4386 1549
rect 4386 1530 4400 1549
rect 4456 1530 4476 1549
rect 4476 1530 4490 1549
rect 4546 1530 4566 1549
rect 4566 1530 4580 1549
rect 4636 1530 4656 1549
rect 4656 1530 4670 1549
rect 4726 1530 4746 1549
rect 4746 1530 4760 1549
rect 4816 1530 4836 1549
rect 4836 1530 4850 1549
rect 4906 1530 4926 1549
rect 4926 1530 4940 1549
rect 4996 1530 5016 1549
rect 5016 1530 5030 1549
rect 5086 1530 5106 1549
rect 5106 1530 5120 1549
rect 5176 1530 5196 1549
rect 5196 1530 5210 1549
rect 5266 1530 5286 1549
rect 5286 1530 5300 1549
rect 5356 1530 5390 1564
rect 5526 1530 5560 1564
rect 5616 1549 5650 1564
rect 5706 1549 5740 1564
rect 5796 1549 5830 1564
rect 5886 1549 5920 1564
rect 5976 1549 6010 1564
rect 6066 1549 6100 1564
rect 6156 1549 6190 1564
rect 6246 1549 6280 1564
rect 6336 1549 6370 1564
rect 6426 1549 6460 1564
rect 6516 1549 6550 1564
rect 6606 1549 6640 1564
rect 5616 1530 5636 1549
rect 5636 1530 5650 1549
rect 5706 1530 5726 1549
rect 5726 1530 5740 1549
rect 5796 1530 5816 1549
rect 5816 1530 5830 1549
rect 5886 1530 5906 1549
rect 5906 1530 5920 1549
rect 5976 1530 5996 1549
rect 5996 1530 6010 1549
rect 6066 1530 6086 1549
rect 6086 1530 6100 1549
rect 6156 1530 6176 1549
rect 6176 1530 6190 1549
rect 6246 1530 6266 1549
rect 6266 1530 6280 1549
rect 6336 1530 6356 1549
rect 6356 1530 6370 1549
rect 6426 1530 6446 1549
rect 6446 1530 6460 1549
rect 6516 1530 6536 1549
rect 6536 1530 6550 1549
rect 6606 1530 6626 1549
rect 6626 1530 6640 1549
rect 6696 1530 6730 1564
rect 6866 1530 6900 1564
rect 6956 1549 6990 1564
rect 7046 1549 7080 1564
rect 7136 1549 7170 1564
rect 7226 1549 7260 1564
rect 7316 1549 7350 1564
rect 7406 1549 7440 1564
rect 7496 1549 7530 1564
rect 7586 1549 7620 1564
rect 7676 1549 7710 1564
rect 7766 1549 7800 1564
rect 7856 1549 7890 1564
rect 7946 1549 7980 1564
rect 6956 1530 6976 1549
rect 6976 1530 6990 1549
rect 7046 1530 7066 1549
rect 7066 1530 7080 1549
rect 7136 1530 7156 1549
rect 7156 1530 7170 1549
rect 7226 1530 7246 1549
rect 7246 1530 7260 1549
rect 7316 1530 7336 1549
rect 7336 1530 7350 1549
rect 7406 1530 7426 1549
rect 7426 1530 7440 1549
rect 7496 1530 7516 1549
rect 7516 1530 7530 1549
rect 7586 1530 7606 1549
rect 7606 1530 7620 1549
rect 7676 1530 7696 1549
rect 7696 1530 7710 1549
rect 7766 1530 7786 1549
rect 7786 1530 7800 1549
rect 7856 1530 7876 1549
rect 7876 1530 7890 1549
rect 7946 1530 7966 1549
rect 7966 1530 7980 1549
rect 8036 1530 8070 1564
rect 8206 1530 8240 1564
rect 8296 1549 8330 1564
rect 8386 1549 8420 1564
rect 8476 1549 8510 1564
rect 8566 1549 8600 1564
rect 8656 1549 8690 1564
rect 8746 1549 8780 1564
rect 8836 1549 8870 1564
rect 8926 1549 8960 1564
rect 9016 1549 9050 1564
rect 9106 1549 9140 1564
rect 9196 1549 9230 1564
rect 9286 1549 9320 1564
rect 8296 1530 8316 1549
rect 8316 1530 8330 1549
rect 8386 1530 8406 1549
rect 8406 1530 8420 1549
rect 8476 1530 8496 1549
rect 8496 1530 8510 1549
rect 8566 1530 8586 1549
rect 8586 1530 8600 1549
rect 8656 1530 8676 1549
rect 8676 1530 8690 1549
rect 8746 1530 8766 1549
rect 8766 1530 8780 1549
rect 8836 1530 8856 1549
rect 8856 1530 8870 1549
rect 8926 1530 8946 1549
rect 8946 1530 8960 1549
rect 9016 1530 9036 1549
rect 9036 1530 9050 1549
rect 9106 1530 9126 1549
rect 9126 1530 9140 1549
rect 9196 1530 9216 1549
rect 9216 1530 9230 1549
rect 9286 1530 9306 1549
rect 9306 1530 9320 1549
rect 9376 1530 9410 1564
rect 9546 1530 9580 1564
rect 9636 1549 9670 1564
rect 9726 1549 9760 1564
rect 9816 1549 9850 1564
rect 9906 1549 9940 1564
rect 9996 1549 10030 1564
rect 10086 1549 10120 1564
rect 10176 1549 10210 1564
rect 10266 1549 10300 1564
rect 10356 1549 10390 1564
rect 10446 1549 10480 1564
rect 10536 1549 10570 1564
rect 10626 1549 10660 1564
rect 9636 1530 9656 1549
rect 9656 1530 9670 1549
rect 9726 1530 9746 1549
rect 9746 1530 9760 1549
rect 9816 1530 9836 1549
rect 9836 1530 9850 1549
rect 9906 1530 9926 1549
rect 9926 1530 9940 1549
rect 9996 1530 10016 1549
rect 10016 1530 10030 1549
rect 10086 1530 10106 1549
rect 10106 1530 10120 1549
rect 10176 1530 10196 1549
rect 10196 1530 10210 1549
rect 10266 1530 10286 1549
rect 10286 1530 10300 1549
rect 10356 1530 10376 1549
rect 10376 1530 10390 1549
rect 10446 1530 10466 1549
rect 10466 1530 10480 1549
rect 10536 1530 10556 1549
rect 10556 1530 10570 1549
rect 10626 1530 10646 1549
rect 10646 1530 10660 1549
rect 10716 1530 10750 1564
rect 330 1370 364 1404
rect 420 1402 454 1404
rect 510 1402 544 1404
rect 600 1402 634 1404
rect 690 1402 724 1404
rect 780 1402 814 1404
rect 870 1402 904 1404
rect 960 1402 994 1404
rect 1050 1402 1084 1404
rect 1140 1402 1174 1404
rect 420 1370 440 1402
rect 440 1370 454 1402
rect 510 1370 530 1402
rect 530 1370 544 1402
rect 600 1370 620 1402
rect 620 1370 634 1402
rect 690 1370 710 1402
rect 710 1370 724 1402
rect 780 1370 800 1402
rect 800 1370 814 1402
rect 870 1370 890 1402
rect 890 1370 904 1402
rect 960 1370 980 1402
rect 980 1370 994 1402
rect 1050 1370 1070 1402
rect 1070 1370 1084 1402
rect 1140 1370 1160 1402
rect 1160 1370 1174 1402
rect 1230 1370 1264 1404
rect 516 1194 538 1200
rect 538 1194 550 1200
rect 616 1194 628 1200
rect 628 1194 650 1200
rect 716 1194 718 1200
rect 718 1194 750 1200
rect 516 1166 550 1194
rect 616 1166 650 1194
rect 716 1166 750 1194
rect 816 1166 850 1200
rect 916 1166 950 1200
rect 1016 1194 1044 1200
rect 1044 1194 1050 1200
rect 1016 1166 1050 1194
rect 516 1066 550 1100
rect 616 1066 650 1100
rect 716 1066 750 1100
rect 816 1066 850 1100
rect 916 1066 950 1100
rect 1016 1066 1050 1100
rect 516 966 550 1000
rect 616 966 650 1000
rect 716 966 750 1000
rect 816 966 850 1000
rect 916 966 950 1000
rect 1016 966 1050 1000
rect 516 868 550 900
rect 616 868 650 900
rect 716 868 750 900
rect 516 866 538 868
rect 538 866 550 868
rect 616 866 628 868
rect 628 866 650 868
rect 716 866 718 868
rect 718 866 750 868
rect 816 866 850 900
rect 916 866 950 900
rect 1016 868 1050 900
rect 1016 866 1044 868
rect 1044 866 1050 868
rect 516 778 550 800
rect 616 778 650 800
rect 716 778 750 800
rect 516 766 538 778
rect 538 766 550 778
rect 616 766 628 778
rect 628 766 650 778
rect 716 766 718 778
rect 718 766 750 778
rect 816 766 850 800
rect 916 766 950 800
rect 1016 778 1050 800
rect 1016 766 1044 778
rect 1044 766 1050 778
rect 516 688 550 700
rect 616 688 650 700
rect 716 688 750 700
rect 516 666 538 688
rect 538 666 550 688
rect 616 666 628 688
rect 628 666 650 688
rect 716 666 718 688
rect 718 666 750 688
rect 816 666 850 700
rect 916 666 950 700
rect 1016 688 1050 700
rect 1016 666 1044 688
rect 1044 666 1050 688
rect 1670 1370 1704 1404
rect 1760 1402 1794 1404
rect 1850 1402 1884 1404
rect 1940 1402 1974 1404
rect 2030 1402 2064 1404
rect 2120 1402 2154 1404
rect 2210 1402 2244 1404
rect 2300 1402 2334 1404
rect 2390 1402 2424 1404
rect 2480 1402 2514 1404
rect 1760 1370 1780 1402
rect 1780 1370 1794 1402
rect 1850 1370 1870 1402
rect 1870 1370 1884 1402
rect 1940 1370 1960 1402
rect 1960 1370 1974 1402
rect 2030 1370 2050 1402
rect 2050 1370 2064 1402
rect 2120 1370 2140 1402
rect 2140 1370 2154 1402
rect 2210 1370 2230 1402
rect 2230 1370 2244 1402
rect 2300 1370 2320 1402
rect 2320 1370 2334 1402
rect 2390 1370 2410 1402
rect 2410 1370 2424 1402
rect 2480 1370 2500 1402
rect 2500 1370 2514 1402
rect 2570 1370 2604 1404
rect 1856 1194 1878 1200
rect 1878 1194 1890 1200
rect 1956 1194 1968 1200
rect 1968 1194 1990 1200
rect 2056 1194 2058 1200
rect 2058 1194 2090 1200
rect 1856 1166 1890 1194
rect 1956 1166 1990 1194
rect 2056 1166 2090 1194
rect 2156 1166 2190 1200
rect 2256 1166 2290 1200
rect 2356 1194 2384 1200
rect 2384 1194 2390 1200
rect 2356 1166 2390 1194
rect 1856 1066 1890 1100
rect 1956 1066 1990 1100
rect 2056 1066 2090 1100
rect 2156 1066 2190 1100
rect 2256 1066 2290 1100
rect 2356 1066 2390 1100
rect 1856 966 1890 1000
rect 1956 966 1990 1000
rect 2056 966 2090 1000
rect 2156 966 2190 1000
rect 2256 966 2290 1000
rect 2356 966 2390 1000
rect 1856 868 1890 900
rect 1956 868 1990 900
rect 2056 868 2090 900
rect 1856 866 1878 868
rect 1878 866 1890 868
rect 1956 866 1968 868
rect 1968 866 1990 868
rect 2056 866 2058 868
rect 2058 866 2090 868
rect 2156 866 2190 900
rect 2256 866 2290 900
rect 2356 868 2390 900
rect 2356 866 2384 868
rect 2384 866 2390 868
rect 1856 778 1890 800
rect 1956 778 1990 800
rect 2056 778 2090 800
rect 1856 766 1878 778
rect 1878 766 1890 778
rect 1956 766 1968 778
rect 1968 766 1990 778
rect 2056 766 2058 778
rect 2058 766 2090 778
rect 2156 766 2190 800
rect 2256 766 2290 800
rect 2356 778 2390 800
rect 2356 766 2384 778
rect 2384 766 2390 778
rect 1856 688 1890 700
rect 1956 688 1990 700
rect 2056 688 2090 700
rect 1856 666 1878 688
rect 1878 666 1890 688
rect 1956 666 1968 688
rect 1968 666 1990 688
rect 2056 666 2058 688
rect 2058 666 2090 688
rect 2156 666 2190 700
rect 2256 666 2290 700
rect 2356 688 2390 700
rect 2356 666 2384 688
rect 2384 666 2390 688
rect 3010 1370 3044 1404
rect 3100 1402 3134 1404
rect 3190 1402 3224 1404
rect 3280 1402 3314 1404
rect 3370 1402 3404 1404
rect 3460 1402 3494 1404
rect 3550 1402 3584 1404
rect 3640 1402 3674 1404
rect 3730 1402 3764 1404
rect 3820 1402 3854 1404
rect 3100 1370 3120 1402
rect 3120 1370 3134 1402
rect 3190 1370 3210 1402
rect 3210 1370 3224 1402
rect 3280 1370 3300 1402
rect 3300 1370 3314 1402
rect 3370 1370 3390 1402
rect 3390 1370 3404 1402
rect 3460 1370 3480 1402
rect 3480 1370 3494 1402
rect 3550 1370 3570 1402
rect 3570 1370 3584 1402
rect 3640 1370 3660 1402
rect 3660 1370 3674 1402
rect 3730 1370 3750 1402
rect 3750 1370 3764 1402
rect 3820 1370 3840 1402
rect 3840 1370 3854 1402
rect 3910 1370 3944 1404
rect 3196 1194 3218 1200
rect 3218 1194 3230 1200
rect 3296 1194 3308 1200
rect 3308 1194 3330 1200
rect 3396 1194 3398 1200
rect 3398 1194 3430 1200
rect 3196 1166 3230 1194
rect 3296 1166 3330 1194
rect 3396 1166 3430 1194
rect 3496 1166 3530 1200
rect 3596 1166 3630 1200
rect 3696 1194 3724 1200
rect 3724 1194 3730 1200
rect 3696 1166 3730 1194
rect 3196 1066 3230 1100
rect 3296 1066 3330 1100
rect 3396 1066 3430 1100
rect 3496 1066 3530 1100
rect 3596 1066 3630 1100
rect 3696 1066 3730 1100
rect 3196 966 3230 1000
rect 3296 966 3330 1000
rect 3396 966 3430 1000
rect 3496 966 3530 1000
rect 3596 966 3630 1000
rect 3696 966 3730 1000
rect 3196 868 3230 900
rect 3296 868 3330 900
rect 3396 868 3430 900
rect 3196 866 3218 868
rect 3218 866 3230 868
rect 3296 866 3308 868
rect 3308 866 3330 868
rect 3396 866 3398 868
rect 3398 866 3430 868
rect 3496 866 3530 900
rect 3596 866 3630 900
rect 3696 868 3730 900
rect 3696 866 3724 868
rect 3724 866 3730 868
rect 3196 778 3230 800
rect 3296 778 3330 800
rect 3396 778 3430 800
rect 3196 766 3218 778
rect 3218 766 3230 778
rect 3296 766 3308 778
rect 3308 766 3330 778
rect 3396 766 3398 778
rect 3398 766 3430 778
rect 3496 766 3530 800
rect 3596 766 3630 800
rect 3696 778 3730 800
rect 3696 766 3724 778
rect 3724 766 3730 778
rect 3196 688 3230 700
rect 3296 688 3330 700
rect 3396 688 3430 700
rect 3196 666 3218 688
rect 3218 666 3230 688
rect 3296 666 3308 688
rect 3308 666 3330 688
rect 3396 666 3398 688
rect 3398 666 3430 688
rect 3496 666 3530 700
rect 3596 666 3630 700
rect 3696 688 3730 700
rect 3696 666 3724 688
rect 3724 666 3730 688
rect 4350 1370 4384 1404
rect 4440 1402 4474 1404
rect 4530 1402 4564 1404
rect 4620 1402 4654 1404
rect 4710 1402 4744 1404
rect 4800 1402 4834 1404
rect 4890 1402 4924 1404
rect 4980 1402 5014 1404
rect 5070 1402 5104 1404
rect 5160 1402 5194 1404
rect 4440 1370 4460 1402
rect 4460 1370 4474 1402
rect 4530 1370 4550 1402
rect 4550 1370 4564 1402
rect 4620 1370 4640 1402
rect 4640 1370 4654 1402
rect 4710 1370 4730 1402
rect 4730 1370 4744 1402
rect 4800 1370 4820 1402
rect 4820 1370 4834 1402
rect 4890 1370 4910 1402
rect 4910 1370 4924 1402
rect 4980 1370 5000 1402
rect 5000 1370 5014 1402
rect 5070 1370 5090 1402
rect 5090 1370 5104 1402
rect 5160 1370 5180 1402
rect 5180 1370 5194 1402
rect 5250 1370 5284 1404
rect 4536 1194 4558 1200
rect 4558 1194 4570 1200
rect 4636 1194 4648 1200
rect 4648 1194 4670 1200
rect 4736 1194 4738 1200
rect 4738 1194 4770 1200
rect 4536 1166 4570 1194
rect 4636 1166 4670 1194
rect 4736 1166 4770 1194
rect 4836 1166 4870 1200
rect 4936 1166 4970 1200
rect 5036 1194 5064 1200
rect 5064 1194 5070 1200
rect 5036 1166 5070 1194
rect 4536 1066 4570 1100
rect 4636 1066 4670 1100
rect 4736 1066 4770 1100
rect 4836 1066 4870 1100
rect 4936 1066 4970 1100
rect 5036 1066 5070 1100
rect 4536 966 4570 1000
rect 4636 966 4670 1000
rect 4736 966 4770 1000
rect 4836 966 4870 1000
rect 4936 966 4970 1000
rect 5036 966 5070 1000
rect 4536 868 4570 900
rect 4636 868 4670 900
rect 4736 868 4770 900
rect 4536 866 4558 868
rect 4558 866 4570 868
rect 4636 866 4648 868
rect 4648 866 4670 868
rect 4736 866 4738 868
rect 4738 866 4770 868
rect 4836 866 4870 900
rect 4936 866 4970 900
rect 5036 868 5070 900
rect 5036 866 5064 868
rect 5064 866 5070 868
rect 4536 778 4570 800
rect 4636 778 4670 800
rect 4736 778 4770 800
rect 4536 766 4558 778
rect 4558 766 4570 778
rect 4636 766 4648 778
rect 4648 766 4670 778
rect 4736 766 4738 778
rect 4738 766 4770 778
rect 4836 766 4870 800
rect 4936 766 4970 800
rect 5036 778 5070 800
rect 5036 766 5064 778
rect 5064 766 5070 778
rect 4536 688 4570 700
rect 4636 688 4670 700
rect 4736 688 4770 700
rect 4536 666 4558 688
rect 4558 666 4570 688
rect 4636 666 4648 688
rect 4648 666 4670 688
rect 4736 666 4738 688
rect 4738 666 4770 688
rect 4836 666 4870 700
rect 4936 666 4970 700
rect 5036 688 5070 700
rect 5036 666 5064 688
rect 5064 666 5070 688
rect 5690 1370 5724 1404
rect 5780 1402 5814 1404
rect 5870 1402 5904 1404
rect 5960 1402 5994 1404
rect 6050 1402 6084 1404
rect 6140 1402 6174 1404
rect 6230 1402 6264 1404
rect 6320 1402 6354 1404
rect 6410 1402 6444 1404
rect 6500 1402 6534 1404
rect 5780 1370 5800 1402
rect 5800 1370 5814 1402
rect 5870 1370 5890 1402
rect 5890 1370 5904 1402
rect 5960 1370 5980 1402
rect 5980 1370 5994 1402
rect 6050 1370 6070 1402
rect 6070 1370 6084 1402
rect 6140 1370 6160 1402
rect 6160 1370 6174 1402
rect 6230 1370 6250 1402
rect 6250 1370 6264 1402
rect 6320 1370 6340 1402
rect 6340 1370 6354 1402
rect 6410 1370 6430 1402
rect 6430 1370 6444 1402
rect 6500 1370 6520 1402
rect 6520 1370 6534 1402
rect 6590 1370 6624 1404
rect 5876 1194 5898 1200
rect 5898 1194 5910 1200
rect 5976 1194 5988 1200
rect 5988 1194 6010 1200
rect 6076 1194 6078 1200
rect 6078 1194 6110 1200
rect 5876 1166 5910 1194
rect 5976 1166 6010 1194
rect 6076 1166 6110 1194
rect 6176 1166 6210 1200
rect 6276 1166 6310 1200
rect 6376 1194 6404 1200
rect 6404 1194 6410 1200
rect 6376 1166 6410 1194
rect 5876 1066 5910 1100
rect 5976 1066 6010 1100
rect 6076 1066 6110 1100
rect 6176 1066 6210 1100
rect 6276 1066 6310 1100
rect 6376 1066 6410 1100
rect 5876 966 5910 1000
rect 5976 966 6010 1000
rect 6076 966 6110 1000
rect 6176 966 6210 1000
rect 6276 966 6310 1000
rect 6376 966 6410 1000
rect 5876 868 5910 900
rect 5976 868 6010 900
rect 6076 868 6110 900
rect 5876 866 5898 868
rect 5898 866 5910 868
rect 5976 866 5988 868
rect 5988 866 6010 868
rect 6076 866 6078 868
rect 6078 866 6110 868
rect 6176 866 6210 900
rect 6276 866 6310 900
rect 6376 868 6410 900
rect 6376 866 6404 868
rect 6404 866 6410 868
rect 5876 778 5910 800
rect 5976 778 6010 800
rect 6076 778 6110 800
rect 5876 766 5898 778
rect 5898 766 5910 778
rect 5976 766 5988 778
rect 5988 766 6010 778
rect 6076 766 6078 778
rect 6078 766 6110 778
rect 6176 766 6210 800
rect 6276 766 6310 800
rect 6376 778 6410 800
rect 6376 766 6404 778
rect 6404 766 6410 778
rect 5876 688 5910 700
rect 5976 688 6010 700
rect 6076 688 6110 700
rect 5876 666 5898 688
rect 5898 666 5910 688
rect 5976 666 5988 688
rect 5988 666 6010 688
rect 6076 666 6078 688
rect 6078 666 6110 688
rect 6176 666 6210 700
rect 6276 666 6310 700
rect 6376 688 6410 700
rect 6376 666 6404 688
rect 6404 666 6410 688
rect 7030 1370 7064 1404
rect 7120 1402 7154 1404
rect 7210 1402 7244 1404
rect 7300 1402 7334 1404
rect 7390 1402 7424 1404
rect 7480 1402 7514 1404
rect 7570 1402 7604 1404
rect 7660 1402 7694 1404
rect 7750 1402 7784 1404
rect 7840 1402 7874 1404
rect 7120 1370 7140 1402
rect 7140 1370 7154 1402
rect 7210 1370 7230 1402
rect 7230 1370 7244 1402
rect 7300 1370 7320 1402
rect 7320 1370 7334 1402
rect 7390 1370 7410 1402
rect 7410 1370 7424 1402
rect 7480 1370 7500 1402
rect 7500 1370 7514 1402
rect 7570 1370 7590 1402
rect 7590 1370 7604 1402
rect 7660 1370 7680 1402
rect 7680 1370 7694 1402
rect 7750 1370 7770 1402
rect 7770 1370 7784 1402
rect 7840 1370 7860 1402
rect 7860 1370 7874 1402
rect 7930 1370 7964 1404
rect 7216 1194 7238 1200
rect 7238 1194 7250 1200
rect 7316 1194 7328 1200
rect 7328 1194 7350 1200
rect 7416 1194 7418 1200
rect 7418 1194 7450 1200
rect 7216 1166 7250 1194
rect 7316 1166 7350 1194
rect 7416 1166 7450 1194
rect 7516 1166 7550 1200
rect 7616 1166 7650 1200
rect 7716 1194 7744 1200
rect 7744 1194 7750 1200
rect 7716 1166 7750 1194
rect 7216 1066 7250 1100
rect 7316 1066 7350 1100
rect 7416 1066 7450 1100
rect 7516 1066 7550 1100
rect 7616 1066 7650 1100
rect 7716 1066 7750 1100
rect 7216 966 7250 1000
rect 7316 966 7350 1000
rect 7416 966 7450 1000
rect 7516 966 7550 1000
rect 7616 966 7650 1000
rect 7716 966 7750 1000
rect 7216 868 7250 900
rect 7316 868 7350 900
rect 7416 868 7450 900
rect 7216 866 7238 868
rect 7238 866 7250 868
rect 7316 866 7328 868
rect 7328 866 7350 868
rect 7416 866 7418 868
rect 7418 866 7450 868
rect 7516 866 7550 900
rect 7616 866 7650 900
rect 7716 868 7750 900
rect 7716 866 7744 868
rect 7744 866 7750 868
rect 7216 778 7250 800
rect 7316 778 7350 800
rect 7416 778 7450 800
rect 7216 766 7238 778
rect 7238 766 7250 778
rect 7316 766 7328 778
rect 7328 766 7350 778
rect 7416 766 7418 778
rect 7418 766 7450 778
rect 7516 766 7550 800
rect 7616 766 7650 800
rect 7716 778 7750 800
rect 7716 766 7744 778
rect 7744 766 7750 778
rect 7216 688 7250 700
rect 7316 688 7350 700
rect 7416 688 7450 700
rect 7216 666 7238 688
rect 7238 666 7250 688
rect 7316 666 7328 688
rect 7328 666 7350 688
rect 7416 666 7418 688
rect 7418 666 7450 688
rect 7516 666 7550 700
rect 7616 666 7650 700
rect 7716 688 7750 700
rect 7716 666 7744 688
rect 7744 666 7750 688
rect 8370 1370 8404 1404
rect 8460 1402 8494 1404
rect 8550 1402 8584 1404
rect 8640 1402 8674 1404
rect 8730 1402 8764 1404
rect 8820 1402 8854 1404
rect 8910 1402 8944 1404
rect 9000 1402 9034 1404
rect 9090 1402 9124 1404
rect 9180 1402 9214 1404
rect 8460 1370 8480 1402
rect 8480 1370 8494 1402
rect 8550 1370 8570 1402
rect 8570 1370 8584 1402
rect 8640 1370 8660 1402
rect 8660 1370 8674 1402
rect 8730 1370 8750 1402
rect 8750 1370 8764 1402
rect 8820 1370 8840 1402
rect 8840 1370 8854 1402
rect 8910 1370 8930 1402
rect 8930 1370 8944 1402
rect 9000 1370 9020 1402
rect 9020 1370 9034 1402
rect 9090 1370 9110 1402
rect 9110 1370 9124 1402
rect 9180 1370 9200 1402
rect 9200 1370 9214 1402
rect 9270 1370 9304 1404
rect 8556 1194 8578 1200
rect 8578 1194 8590 1200
rect 8656 1194 8668 1200
rect 8668 1194 8690 1200
rect 8756 1194 8758 1200
rect 8758 1194 8790 1200
rect 8556 1166 8590 1194
rect 8656 1166 8690 1194
rect 8756 1166 8790 1194
rect 8856 1166 8890 1200
rect 8956 1166 8990 1200
rect 9056 1194 9084 1200
rect 9084 1194 9090 1200
rect 9056 1166 9090 1194
rect 8556 1066 8590 1100
rect 8656 1066 8690 1100
rect 8756 1066 8790 1100
rect 8856 1066 8890 1100
rect 8956 1066 8990 1100
rect 9056 1066 9090 1100
rect 8556 966 8590 1000
rect 8656 966 8690 1000
rect 8756 966 8790 1000
rect 8856 966 8890 1000
rect 8956 966 8990 1000
rect 9056 966 9090 1000
rect 8556 868 8590 900
rect 8656 868 8690 900
rect 8756 868 8790 900
rect 8556 866 8578 868
rect 8578 866 8590 868
rect 8656 866 8668 868
rect 8668 866 8690 868
rect 8756 866 8758 868
rect 8758 866 8790 868
rect 8856 866 8890 900
rect 8956 866 8990 900
rect 9056 868 9090 900
rect 9056 866 9084 868
rect 9084 866 9090 868
rect 8556 778 8590 800
rect 8656 778 8690 800
rect 8756 778 8790 800
rect 8556 766 8578 778
rect 8578 766 8590 778
rect 8656 766 8668 778
rect 8668 766 8690 778
rect 8756 766 8758 778
rect 8758 766 8790 778
rect 8856 766 8890 800
rect 8956 766 8990 800
rect 9056 778 9090 800
rect 9056 766 9084 778
rect 9084 766 9090 778
rect 8556 688 8590 700
rect 8656 688 8690 700
rect 8756 688 8790 700
rect 8556 666 8578 688
rect 8578 666 8590 688
rect 8656 666 8668 688
rect 8668 666 8690 688
rect 8756 666 8758 688
rect 8758 666 8790 688
rect 8856 666 8890 700
rect 8956 666 8990 700
rect 9056 688 9090 700
rect 9056 666 9084 688
rect 9084 666 9090 688
rect 9710 1370 9744 1404
rect 9800 1402 9834 1404
rect 9890 1402 9924 1404
rect 9980 1402 10014 1404
rect 10070 1402 10104 1404
rect 10160 1402 10194 1404
rect 10250 1402 10284 1404
rect 10340 1402 10374 1404
rect 10430 1402 10464 1404
rect 10520 1402 10554 1404
rect 9800 1370 9820 1402
rect 9820 1370 9834 1402
rect 9890 1370 9910 1402
rect 9910 1370 9924 1402
rect 9980 1370 10000 1402
rect 10000 1370 10014 1402
rect 10070 1370 10090 1402
rect 10090 1370 10104 1402
rect 10160 1370 10180 1402
rect 10180 1370 10194 1402
rect 10250 1370 10270 1402
rect 10270 1370 10284 1402
rect 10340 1370 10360 1402
rect 10360 1370 10374 1402
rect 10430 1370 10450 1402
rect 10450 1370 10464 1402
rect 10520 1370 10540 1402
rect 10540 1370 10554 1402
rect 10610 1370 10644 1404
rect 9896 1194 9918 1200
rect 9918 1194 9930 1200
rect 9996 1194 10008 1200
rect 10008 1194 10030 1200
rect 10096 1194 10098 1200
rect 10098 1194 10130 1200
rect 9896 1166 9930 1194
rect 9996 1166 10030 1194
rect 10096 1166 10130 1194
rect 10196 1166 10230 1200
rect 10296 1166 10330 1200
rect 10396 1194 10424 1200
rect 10424 1194 10430 1200
rect 10396 1166 10430 1194
rect 9896 1066 9930 1100
rect 9996 1066 10030 1100
rect 10096 1066 10130 1100
rect 10196 1066 10230 1100
rect 10296 1066 10330 1100
rect 10396 1066 10430 1100
rect 9896 966 9930 1000
rect 9996 966 10030 1000
rect 10096 966 10130 1000
rect 10196 966 10230 1000
rect 10296 966 10330 1000
rect 10396 966 10430 1000
rect 9896 868 9930 900
rect 9996 868 10030 900
rect 10096 868 10130 900
rect 9896 866 9918 868
rect 9918 866 9930 868
rect 9996 866 10008 868
rect 10008 866 10030 868
rect 10096 866 10098 868
rect 10098 866 10130 868
rect 10196 866 10230 900
rect 10296 866 10330 900
rect 10396 868 10430 900
rect 10396 866 10424 868
rect 10424 866 10430 868
rect 9896 778 9930 800
rect 9996 778 10030 800
rect 10096 778 10130 800
rect 9896 766 9918 778
rect 9918 766 9930 778
rect 9996 766 10008 778
rect 10008 766 10030 778
rect 10096 766 10098 778
rect 10098 766 10130 778
rect 10196 766 10230 800
rect 10296 766 10330 800
rect 10396 778 10430 800
rect 10396 766 10424 778
rect 10424 766 10430 778
rect 9896 688 9930 700
rect 9996 688 10030 700
rect 10096 688 10130 700
rect 9896 666 9918 688
rect 9918 666 9930 688
rect 9996 666 10008 688
rect 10008 666 10030 688
rect 10096 666 10098 688
rect 10098 666 10130 688
rect 10196 666 10230 700
rect 10296 666 10330 700
rect 10396 688 10430 700
rect 10396 666 10424 688
rect 10424 666 10430 688
rect 303 -17 337 17
rect 503 -17 537 17
rect 703 -17 737 17
rect 903 -17 937 17
rect 1103 -17 1137 17
rect 1303 -17 1337 17
rect 1503 -17 1537 17
rect 1703 -17 1737 17
rect 1903 -17 1937 17
rect 2103 -17 2137 17
rect 2303 -17 2337 17
rect 2503 -17 2537 17
rect 2703 -17 2737 17
rect 2903 -17 2937 17
rect 3103 -17 3137 17
rect 3303 -17 3337 17
rect 3503 -17 3537 17
rect 3703 -17 3737 17
rect 3903 -17 3937 17
rect 4103 -17 4137 17
rect 4303 -17 4337 17
rect 4503 -17 4537 17
rect 4703 -17 4737 17
rect 4903 -17 4937 17
rect 5103 -17 5137 17
rect 5303 -17 5337 17
rect 5503 -17 5537 17
rect 5703 -17 5737 17
rect 5903 -17 5937 17
rect 6103 -17 6137 17
rect 6303 -17 6337 17
rect 6503 -17 6537 17
rect 6703 -17 6737 17
rect 6903 -17 6937 17
rect 7103 -17 7137 17
rect 7303 -17 7337 17
rect 7503 -17 7537 17
rect 7703 -17 7737 17
rect 7903 -17 7937 17
rect 8103 -17 8137 17
rect 8303 -17 8337 17
rect 8503 -17 8537 17
rect 8703 -17 8737 17
rect 8903 -17 8937 17
rect 9103 -17 9137 17
rect 9303 -17 9337 17
rect 9503 -17 9537 17
rect 9703 -17 9737 17
rect 9903 -17 9937 17
rect 10103 -17 10137 17
rect 10303 -17 10337 17
rect 10503 -17 10537 17
rect 10703 -17 10737 17
<< metal1 >>
rect 120 1897 10840 1940
rect 120 1863 303 1897
rect 337 1863 503 1897
rect 537 1863 703 1897
rect 737 1863 903 1897
rect 937 1863 1103 1897
rect 1137 1863 1303 1897
rect 1337 1863 1503 1897
rect 1537 1863 1703 1897
rect 1737 1863 1903 1897
rect 1937 1863 2103 1897
rect 2137 1863 2303 1897
rect 2337 1863 2503 1897
rect 2537 1863 2703 1897
rect 2737 1863 2903 1897
rect 2937 1863 3103 1897
rect 3137 1863 3303 1897
rect 3337 1863 3503 1897
rect 3537 1863 3703 1897
rect 3737 1863 3903 1897
rect 3937 1863 4103 1897
rect 4137 1863 4303 1897
rect 4337 1863 4503 1897
rect 4537 1863 4703 1897
rect 4737 1863 4903 1897
rect 4937 1863 5103 1897
rect 5137 1863 5303 1897
rect 5337 1863 5503 1897
rect 5537 1863 5703 1897
rect 5737 1863 5903 1897
rect 5937 1863 6103 1897
rect 6137 1863 6303 1897
rect 6337 1863 6503 1897
rect 6537 1863 6703 1897
rect 6737 1863 6903 1897
rect 6937 1863 7103 1897
rect 7137 1863 7303 1897
rect 7337 1863 7503 1897
rect 7537 1863 7703 1897
rect 7737 1863 7903 1897
rect 7937 1863 8103 1897
rect 8137 1863 8303 1897
rect 8337 1863 8503 1897
rect 8537 1863 8703 1897
rect 8737 1863 8903 1897
rect 8937 1863 9103 1897
rect 9137 1863 9303 1897
rect 9337 1863 9503 1897
rect 9537 1863 9703 1897
rect 9737 1863 9903 1897
rect 9937 1863 10103 1897
rect 10137 1863 10303 1897
rect 10337 1863 10503 1897
rect 10537 1863 10703 1897
rect 10737 1863 10840 1897
rect 120 1820 10840 1863
rect 146 1564 10814 1570
rect 146 1530 166 1564
rect 200 1530 256 1564
rect 290 1530 346 1564
rect 380 1530 436 1564
rect 470 1530 526 1564
rect 560 1530 616 1564
rect 650 1530 706 1564
rect 740 1530 796 1564
rect 830 1530 886 1564
rect 920 1530 976 1564
rect 1010 1530 1066 1564
rect 1100 1530 1156 1564
rect 1190 1530 1246 1564
rect 1280 1530 1336 1564
rect 1370 1530 1506 1564
rect 1540 1530 1596 1564
rect 1630 1530 1686 1564
rect 1720 1530 1776 1564
rect 1810 1530 1866 1564
rect 1900 1530 1956 1564
rect 1990 1530 2046 1564
rect 2080 1530 2136 1564
rect 2170 1530 2226 1564
rect 2260 1530 2316 1564
rect 2350 1530 2406 1564
rect 2440 1530 2496 1564
rect 2530 1530 2586 1564
rect 2620 1530 2676 1564
rect 2710 1530 2846 1564
rect 2880 1530 2936 1564
rect 2970 1530 3026 1564
rect 3060 1530 3116 1564
rect 3150 1530 3206 1564
rect 3240 1530 3296 1564
rect 3330 1530 3386 1564
rect 3420 1530 3476 1564
rect 3510 1530 3566 1564
rect 3600 1530 3656 1564
rect 3690 1530 3746 1564
rect 3780 1530 3836 1564
rect 3870 1530 3926 1564
rect 3960 1530 4016 1564
rect 4050 1530 4186 1564
rect 4220 1530 4276 1564
rect 4310 1530 4366 1564
rect 4400 1530 4456 1564
rect 4490 1530 4546 1564
rect 4580 1530 4636 1564
rect 4670 1530 4726 1564
rect 4760 1530 4816 1564
rect 4850 1530 4906 1564
rect 4940 1530 4996 1564
rect 5030 1530 5086 1564
rect 5120 1530 5176 1564
rect 5210 1530 5266 1564
rect 5300 1530 5356 1564
rect 5390 1530 5526 1564
rect 5560 1530 5616 1564
rect 5650 1530 5706 1564
rect 5740 1530 5796 1564
rect 5830 1530 5886 1564
rect 5920 1530 5976 1564
rect 6010 1530 6066 1564
rect 6100 1530 6156 1564
rect 6190 1530 6246 1564
rect 6280 1530 6336 1564
rect 6370 1530 6426 1564
rect 6460 1530 6516 1564
rect 6550 1530 6606 1564
rect 6640 1530 6696 1564
rect 6730 1530 6866 1564
rect 6900 1530 6956 1564
rect 6990 1530 7046 1564
rect 7080 1530 7136 1564
rect 7170 1530 7226 1564
rect 7260 1530 7316 1564
rect 7350 1530 7406 1564
rect 7440 1530 7496 1564
rect 7530 1530 7586 1564
rect 7620 1530 7676 1564
rect 7710 1530 7766 1564
rect 7800 1530 7856 1564
rect 7890 1530 7946 1564
rect 7980 1530 8036 1564
rect 8070 1530 8206 1564
rect 8240 1530 8296 1564
rect 8330 1530 8386 1564
rect 8420 1530 8476 1564
rect 8510 1530 8566 1564
rect 8600 1530 8656 1564
rect 8690 1530 8746 1564
rect 8780 1530 8836 1564
rect 8870 1530 8926 1564
rect 8960 1530 9016 1564
rect 9050 1530 9106 1564
rect 9140 1530 9196 1564
rect 9230 1530 9286 1564
rect 9320 1530 9376 1564
rect 9410 1530 9546 1564
rect 9580 1530 9636 1564
rect 9670 1530 9726 1564
rect 9760 1530 9816 1564
rect 9850 1530 9906 1564
rect 9940 1530 9996 1564
rect 10030 1530 10086 1564
rect 10120 1530 10176 1564
rect 10210 1530 10266 1564
rect 10300 1530 10356 1564
rect 10390 1530 10446 1564
rect 10480 1530 10536 1564
rect 10570 1530 10626 1564
rect 10660 1530 10716 1564
rect 10750 1530 10814 1564
rect 146 1500 10814 1530
rect 310 1404 10650 1420
rect 310 1370 330 1404
rect 364 1370 420 1404
rect 454 1370 510 1404
rect 544 1370 600 1404
rect 634 1370 690 1404
rect 724 1370 780 1404
rect 814 1370 870 1404
rect 904 1370 960 1404
rect 994 1370 1050 1404
rect 1084 1370 1140 1404
rect 1174 1370 1230 1404
rect 1264 1370 1670 1404
rect 1704 1370 1760 1404
rect 1794 1370 1850 1404
rect 1884 1370 1940 1404
rect 1974 1370 2030 1404
rect 2064 1370 2120 1404
rect 2154 1370 2210 1404
rect 2244 1370 2300 1404
rect 2334 1370 2390 1404
rect 2424 1370 2480 1404
rect 2514 1370 2570 1404
rect 2604 1370 3010 1404
rect 3044 1370 3100 1404
rect 3134 1370 3190 1404
rect 3224 1370 3280 1404
rect 3314 1370 3370 1404
rect 3404 1370 3460 1404
rect 3494 1370 3550 1404
rect 3584 1370 3640 1404
rect 3674 1370 3730 1404
rect 3764 1370 3820 1404
rect 3854 1370 3910 1404
rect 3944 1370 4350 1404
rect 4384 1370 4440 1404
rect 4474 1370 4530 1404
rect 4564 1370 4620 1404
rect 4654 1370 4710 1404
rect 4744 1370 4800 1404
rect 4834 1370 4890 1404
rect 4924 1370 4980 1404
rect 5014 1370 5070 1404
rect 5104 1370 5160 1404
rect 5194 1370 5250 1404
rect 5284 1370 5690 1404
rect 5724 1370 5780 1404
rect 5814 1370 5870 1404
rect 5904 1370 5960 1404
rect 5994 1370 6050 1404
rect 6084 1370 6140 1404
rect 6174 1370 6230 1404
rect 6264 1370 6320 1404
rect 6354 1370 6410 1404
rect 6444 1370 6500 1404
rect 6534 1370 6590 1404
rect 6624 1370 7030 1404
rect 7064 1370 7120 1404
rect 7154 1370 7210 1404
rect 7244 1370 7300 1404
rect 7334 1370 7390 1404
rect 7424 1370 7480 1404
rect 7514 1370 7570 1404
rect 7604 1370 7660 1404
rect 7694 1370 7750 1404
rect 7784 1370 7840 1404
rect 7874 1370 7930 1404
rect 7964 1370 8370 1404
rect 8404 1370 8460 1404
rect 8494 1370 8550 1404
rect 8584 1370 8640 1404
rect 8674 1370 8730 1404
rect 8764 1370 8820 1404
rect 8854 1370 8910 1404
rect 8944 1370 9000 1404
rect 9034 1370 9090 1404
rect 9124 1370 9180 1404
rect 9214 1370 9270 1404
rect 9304 1370 9710 1404
rect 9744 1370 9800 1404
rect 9834 1370 9890 1404
rect 9924 1370 9980 1404
rect 10014 1370 10070 1404
rect 10104 1370 10160 1404
rect 10194 1370 10250 1404
rect 10284 1370 10340 1404
rect 10374 1370 10430 1404
rect 10464 1370 10520 1404
rect 10554 1370 10610 1404
rect 10644 1370 10650 1404
rect 310 1350 10650 1370
rect 484 1200 10476 1246
rect 484 1166 516 1200
rect 550 1166 616 1200
rect 650 1166 716 1200
rect 750 1166 816 1200
rect 850 1166 916 1200
rect 950 1166 1016 1200
rect 1050 1166 1856 1200
rect 1890 1166 1956 1200
rect 1990 1166 2056 1200
rect 2090 1166 2156 1200
rect 2190 1166 2256 1200
rect 2290 1166 2356 1200
rect 2390 1166 3196 1200
rect 3230 1166 3296 1200
rect 3330 1166 3396 1200
rect 3430 1166 3496 1200
rect 3530 1166 3596 1200
rect 3630 1166 3696 1200
rect 3730 1166 4536 1200
rect 4570 1166 4636 1200
rect 4670 1166 4736 1200
rect 4770 1166 4836 1200
rect 4870 1166 4936 1200
rect 4970 1166 5036 1200
rect 5070 1166 5876 1200
rect 5910 1166 5976 1200
rect 6010 1166 6076 1200
rect 6110 1166 6176 1200
rect 6210 1166 6276 1200
rect 6310 1166 6376 1200
rect 6410 1166 7216 1200
rect 7250 1166 7316 1200
rect 7350 1166 7416 1200
rect 7450 1166 7516 1200
rect 7550 1166 7616 1200
rect 7650 1166 7716 1200
rect 7750 1166 8556 1200
rect 8590 1166 8656 1200
rect 8690 1166 8756 1200
rect 8790 1166 8856 1200
rect 8890 1166 8956 1200
rect 8990 1166 9056 1200
rect 9090 1166 9896 1200
rect 9930 1166 9996 1200
rect 10030 1166 10096 1200
rect 10130 1166 10196 1200
rect 10230 1166 10296 1200
rect 10330 1166 10396 1200
rect 10430 1166 10476 1200
rect 484 1100 10476 1166
rect 484 1066 516 1100
rect 550 1066 616 1100
rect 650 1066 716 1100
rect 750 1066 816 1100
rect 850 1066 916 1100
rect 950 1066 1016 1100
rect 1050 1066 1856 1100
rect 1890 1066 1956 1100
rect 1990 1066 2056 1100
rect 2090 1066 2156 1100
rect 2190 1066 2256 1100
rect 2290 1066 2356 1100
rect 2390 1066 3196 1100
rect 3230 1066 3296 1100
rect 3330 1066 3396 1100
rect 3430 1066 3496 1100
rect 3530 1066 3596 1100
rect 3630 1066 3696 1100
rect 3730 1066 4536 1100
rect 4570 1066 4636 1100
rect 4670 1066 4736 1100
rect 4770 1066 4836 1100
rect 4870 1066 4936 1100
rect 4970 1066 5036 1100
rect 5070 1066 5876 1100
rect 5910 1066 5976 1100
rect 6010 1066 6076 1100
rect 6110 1066 6176 1100
rect 6210 1066 6276 1100
rect 6310 1066 6376 1100
rect 6410 1066 7216 1100
rect 7250 1066 7316 1100
rect 7350 1066 7416 1100
rect 7450 1066 7516 1100
rect 7550 1066 7616 1100
rect 7650 1066 7716 1100
rect 7750 1066 8556 1100
rect 8590 1066 8656 1100
rect 8690 1066 8756 1100
rect 8790 1066 8856 1100
rect 8890 1066 8956 1100
rect 8990 1066 9056 1100
rect 9090 1066 9896 1100
rect 9930 1066 9996 1100
rect 10030 1066 10096 1100
rect 10130 1066 10196 1100
rect 10230 1066 10296 1100
rect 10330 1066 10396 1100
rect 10430 1066 10476 1100
rect 484 1000 10476 1066
rect 484 966 516 1000
rect 550 966 616 1000
rect 650 966 716 1000
rect 750 966 816 1000
rect 850 966 916 1000
rect 950 966 1016 1000
rect 1050 966 1856 1000
rect 1890 966 1956 1000
rect 1990 966 2056 1000
rect 2090 966 2156 1000
rect 2190 966 2256 1000
rect 2290 966 2356 1000
rect 2390 966 3196 1000
rect 3230 966 3296 1000
rect 3330 966 3396 1000
rect 3430 966 3496 1000
rect 3530 966 3596 1000
rect 3630 966 3696 1000
rect 3730 966 4536 1000
rect 4570 966 4636 1000
rect 4670 966 4736 1000
rect 4770 966 4836 1000
rect 4870 966 4936 1000
rect 4970 966 5036 1000
rect 5070 966 5876 1000
rect 5910 966 5976 1000
rect 6010 966 6076 1000
rect 6110 966 6176 1000
rect 6210 966 6276 1000
rect 6310 966 6376 1000
rect 6410 966 7216 1000
rect 7250 966 7316 1000
rect 7350 966 7416 1000
rect 7450 966 7516 1000
rect 7550 966 7616 1000
rect 7650 966 7716 1000
rect 7750 966 8556 1000
rect 8590 966 8656 1000
rect 8690 966 8756 1000
rect 8790 966 8856 1000
rect 8890 966 8956 1000
rect 8990 966 9056 1000
rect 9090 966 9896 1000
rect 9930 966 9996 1000
rect 10030 966 10096 1000
rect 10130 966 10196 1000
rect 10230 966 10296 1000
rect 10330 966 10396 1000
rect 10430 966 10476 1000
rect 484 900 10476 966
rect 484 866 516 900
rect 550 866 616 900
rect 650 866 716 900
rect 750 866 816 900
rect 850 866 916 900
rect 950 866 1016 900
rect 1050 866 1856 900
rect 1890 866 1956 900
rect 1990 866 2056 900
rect 2090 866 2156 900
rect 2190 866 2256 900
rect 2290 866 2356 900
rect 2390 866 3196 900
rect 3230 866 3296 900
rect 3330 866 3396 900
rect 3430 866 3496 900
rect 3530 866 3596 900
rect 3630 866 3696 900
rect 3730 866 4536 900
rect 4570 866 4636 900
rect 4670 866 4736 900
rect 4770 866 4836 900
rect 4870 866 4936 900
rect 4970 866 5036 900
rect 5070 866 5876 900
rect 5910 866 5976 900
rect 6010 866 6076 900
rect 6110 866 6176 900
rect 6210 866 6276 900
rect 6310 866 6376 900
rect 6410 866 7216 900
rect 7250 866 7316 900
rect 7350 866 7416 900
rect 7450 866 7516 900
rect 7550 866 7616 900
rect 7650 866 7716 900
rect 7750 866 8556 900
rect 8590 866 8656 900
rect 8690 866 8756 900
rect 8790 866 8856 900
rect 8890 866 8956 900
rect 8990 866 9056 900
rect 9090 866 9896 900
rect 9930 866 9996 900
rect 10030 866 10096 900
rect 10130 866 10196 900
rect 10230 866 10296 900
rect 10330 866 10396 900
rect 10430 866 10476 900
rect 484 800 10476 866
rect 484 766 516 800
rect 550 766 616 800
rect 650 766 716 800
rect 750 766 816 800
rect 850 766 916 800
rect 950 766 1016 800
rect 1050 766 1856 800
rect 1890 766 1956 800
rect 1990 766 2056 800
rect 2090 766 2156 800
rect 2190 766 2256 800
rect 2290 766 2356 800
rect 2390 766 3196 800
rect 3230 766 3296 800
rect 3330 766 3396 800
rect 3430 766 3496 800
rect 3530 766 3596 800
rect 3630 766 3696 800
rect 3730 766 4536 800
rect 4570 766 4636 800
rect 4670 766 4736 800
rect 4770 766 4836 800
rect 4870 766 4936 800
rect 4970 766 5036 800
rect 5070 766 5876 800
rect 5910 766 5976 800
rect 6010 766 6076 800
rect 6110 766 6176 800
rect 6210 766 6276 800
rect 6310 766 6376 800
rect 6410 766 7216 800
rect 7250 766 7316 800
rect 7350 766 7416 800
rect 7450 766 7516 800
rect 7550 766 7616 800
rect 7650 766 7716 800
rect 7750 766 8556 800
rect 8590 766 8656 800
rect 8690 766 8756 800
rect 8790 766 8856 800
rect 8890 766 8956 800
rect 8990 766 9056 800
rect 9090 766 9896 800
rect 9930 766 9996 800
rect 10030 766 10096 800
rect 10130 766 10196 800
rect 10230 766 10296 800
rect 10330 766 10396 800
rect 10430 766 10476 800
rect 484 700 10476 766
rect 484 666 516 700
rect 550 666 616 700
rect 650 666 716 700
rect 750 666 816 700
rect 850 666 916 700
rect 950 666 1016 700
rect 1050 666 1856 700
rect 1890 666 1956 700
rect 1990 666 2056 700
rect 2090 666 2156 700
rect 2190 666 2256 700
rect 2290 666 2356 700
rect 2390 666 3196 700
rect 3230 666 3296 700
rect 3330 666 3396 700
rect 3430 666 3496 700
rect 3530 666 3596 700
rect 3630 666 3696 700
rect 3730 666 4536 700
rect 4570 666 4636 700
rect 4670 666 4736 700
rect 4770 666 4836 700
rect 4870 666 4936 700
rect 4970 666 5036 700
rect 5070 666 5876 700
rect 5910 666 5976 700
rect 6010 666 6076 700
rect 6110 666 6176 700
rect 6210 666 6276 700
rect 6310 666 6376 700
rect 6410 666 7216 700
rect 7250 666 7316 700
rect 7350 666 7416 700
rect 7450 666 7516 700
rect 7550 666 7616 700
rect 7650 666 7716 700
rect 7750 666 8556 700
rect 8590 666 8656 700
rect 8690 666 8756 700
rect 8790 666 8856 700
rect 8890 666 8956 700
rect 8990 666 9056 700
rect 9090 666 9896 700
rect 9930 666 9996 700
rect 10030 666 10096 700
rect 10130 666 10196 700
rect 10230 666 10296 700
rect 10330 666 10396 700
rect 10430 666 10476 700
rect 484 634 10476 666
rect 120 17 10840 60
rect 120 -17 303 17
rect 337 -17 503 17
rect 537 -17 703 17
rect 737 -17 903 17
rect 937 -17 1103 17
rect 1137 -17 1303 17
rect 1337 -17 1503 17
rect 1537 -17 1703 17
rect 1737 -17 1903 17
rect 1937 -17 2103 17
rect 2137 -17 2303 17
rect 2337 -17 2503 17
rect 2537 -17 2703 17
rect 2737 -17 2903 17
rect 2937 -17 3103 17
rect 3137 -17 3303 17
rect 3337 -17 3503 17
rect 3537 -17 3703 17
rect 3737 -17 3903 17
rect 3937 -17 4103 17
rect 4137 -17 4303 17
rect 4337 -17 4503 17
rect 4537 -17 4703 17
rect 4737 -17 4903 17
rect 4937 -17 5103 17
rect 5137 -17 5303 17
rect 5337 -17 5503 17
rect 5537 -17 5703 17
rect 5737 -17 5903 17
rect 5937 -17 6103 17
rect 6137 -17 6303 17
rect 6337 -17 6503 17
rect 6537 -17 6703 17
rect 6737 -17 6903 17
rect 6937 -17 7103 17
rect 7137 -17 7303 17
rect 7337 -17 7503 17
rect 7537 -17 7703 17
rect 7737 -17 7903 17
rect 7937 -17 8103 17
rect 8137 -17 8303 17
rect 8337 -17 8503 17
rect 8537 -17 8703 17
rect 8737 -17 8903 17
rect 8937 -17 9103 17
rect 9137 -17 9303 17
rect 9337 -17 9503 17
rect 9537 -17 9703 17
rect 9737 -17 9903 17
rect 9937 -17 10103 17
rect 10137 -17 10303 17
rect 10337 -17 10503 17
rect 10537 -17 10703 17
rect 10737 -17 10840 17
rect 120 -60 10840 -17
<< labels >>
flabel locali s 10054 896 10302 1000 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
port 1 nsew
flabel locali s 10113 1522 10214 1571 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
port 2 nsew
flabel locali s 10090 1372 10208 1412 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
port 3 nsew
flabel locali s 8714 896 8962 1000 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
port 4 nsew
flabel locali s 8773 1522 8874 1571 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
port 5 nsew
flabel locali s 8750 1372 8868 1412 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
port 6 nsew
flabel locali s 7374 896 7622 1000 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
port 7 nsew
flabel locali s 7433 1522 7534 1571 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
port 8 nsew
flabel locali s 7410 1372 7528 1412 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
port 9 nsew
flabel locali s 6034 896 6282 1000 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
port 10 nsew
flabel locali s 6093 1522 6194 1571 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
port 11 nsew
flabel locali s 6070 1372 6188 1412 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
port 12 nsew
flabel locali s 4694 896 4942 1000 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
port 13 nsew
flabel locali s 4753 1522 4854 1571 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
port 14 nsew
flabel locali s 4730 1372 4848 1412 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
port 15 nsew
flabel locali s 3354 896 3602 1000 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
port 16 nsew
flabel locali s 3413 1522 3514 1571 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
port 17 nsew
flabel locali s 3390 1372 3508 1412 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
port 18 nsew
flabel locali s 2014 896 2262 1000 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
port 19 nsew
flabel locali s 2073 1522 2174 1571 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
port 20 nsew
flabel locali s 2050 1372 2168 1412 0 FreeSans 625 0 0 0 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
port 21 nsew
flabel locali s 674 896 922 1000 0 FreeSans 625 0 0 0 xm1/Emitter
port 22 nsew
flabel locali s 733 1522 834 1571 0 FreeSans 625 0 0 0 xm1/Collector
port 23 nsew
flabel locali s 710 1372 828 1412 0 FreeSans 625 0 0 0 xm1/Base
port 24 nsew
flabel metal1 s 660 1010 900 1140 1 FreeSans 750 0 0 0 Emitter
port 25 nsew
flabel metal1 s 310 1372 550 1412 1 FreeSans 750 0 0 0 Base
port 26 nsew
flabel metal1 s 146 1524 386 1564 1 FreeSans 750 0 0 0 Collector
port 27 nsew
flabel metal1 s 120 1850 180 1910 1 FreeSans 1250 0 0 0 VPWR
port 28 nsew
flabel metal1 s 120 -30 180 30 1 FreeSans 1250 0 0 0 VGND
port 29 nsew
<< properties >>
string FIXED_BBOX 0 0 10960 1880
<< end >>
