magic
tech sky130A
magscale 1 2
timestamp 1655770899
<< pwell >>
rect 134 1426 4420 1500
rect 134 574 4424 1426
rect 134 226 4420 574
rect 132 54 4420 226
rect 134 -52 4420 54
<< nmoslvt >>
rect 276 600 676 1400
rect 734 600 1134 1400
rect 1192 600 1592 1400
rect 1650 600 2050 1400
rect 2108 600 2508 1400
rect 2566 600 2966 1400
rect 3024 600 3424 1400
rect 3482 600 3882 1400
rect 3940 600 4340 1400
<< ndiff >>
rect 218 1357 276 1400
rect 218 1323 230 1357
rect 264 1323 276 1357
rect 218 1289 276 1323
rect 218 1255 230 1289
rect 264 1255 276 1289
rect 218 1221 276 1255
rect 218 1187 230 1221
rect 264 1187 276 1221
rect 218 1153 276 1187
rect 218 1119 230 1153
rect 264 1119 276 1153
rect 218 1085 276 1119
rect 218 1051 230 1085
rect 264 1051 276 1085
rect 218 1017 276 1051
rect 218 983 230 1017
rect 264 983 276 1017
rect 218 949 276 983
rect 218 915 230 949
rect 264 915 276 949
rect 218 881 276 915
rect 218 847 230 881
rect 264 847 276 881
rect 218 813 276 847
rect 218 779 230 813
rect 264 779 276 813
rect 218 745 276 779
rect 218 711 230 745
rect 264 711 276 745
rect 218 677 276 711
rect 218 643 230 677
rect 264 643 276 677
rect 218 600 276 643
rect 676 1357 734 1400
rect 676 1323 688 1357
rect 722 1323 734 1357
rect 676 1289 734 1323
rect 676 1255 688 1289
rect 722 1255 734 1289
rect 676 1221 734 1255
rect 676 1187 688 1221
rect 722 1187 734 1221
rect 676 1153 734 1187
rect 676 1119 688 1153
rect 722 1119 734 1153
rect 676 1085 734 1119
rect 676 1051 688 1085
rect 722 1051 734 1085
rect 676 1017 734 1051
rect 676 983 688 1017
rect 722 983 734 1017
rect 676 949 734 983
rect 676 915 688 949
rect 722 915 734 949
rect 676 881 734 915
rect 676 847 688 881
rect 722 847 734 881
rect 676 813 734 847
rect 676 779 688 813
rect 722 779 734 813
rect 676 745 734 779
rect 676 711 688 745
rect 722 711 734 745
rect 676 677 734 711
rect 676 643 688 677
rect 722 643 734 677
rect 676 600 734 643
rect 1134 1357 1192 1400
rect 1134 1323 1146 1357
rect 1180 1323 1192 1357
rect 1134 1289 1192 1323
rect 1134 1255 1146 1289
rect 1180 1255 1192 1289
rect 1134 1221 1192 1255
rect 1134 1187 1146 1221
rect 1180 1187 1192 1221
rect 1134 1153 1192 1187
rect 1134 1119 1146 1153
rect 1180 1119 1192 1153
rect 1134 1085 1192 1119
rect 1134 1051 1146 1085
rect 1180 1051 1192 1085
rect 1134 1017 1192 1051
rect 1134 983 1146 1017
rect 1180 983 1192 1017
rect 1134 949 1192 983
rect 1134 915 1146 949
rect 1180 915 1192 949
rect 1134 881 1192 915
rect 1134 847 1146 881
rect 1180 847 1192 881
rect 1134 813 1192 847
rect 1134 779 1146 813
rect 1180 779 1192 813
rect 1134 745 1192 779
rect 1134 711 1146 745
rect 1180 711 1192 745
rect 1134 677 1192 711
rect 1134 643 1146 677
rect 1180 643 1192 677
rect 1134 600 1192 643
rect 1592 1357 1650 1400
rect 1592 1323 1604 1357
rect 1638 1323 1650 1357
rect 1592 1289 1650 1323
rect 1592 1255 1604 1289
rect 1638 1255 1650 1289
rect 1592 1221 1650 1255
rect 1592 1187 1604 1221
rect 1638 1187 1650 1221
rect 1592 1153 1650 1187
rect 1592 1119 1604 1153
rect 1638 1119 1650 1153
rect 1592 1085 1650 1119
rect 1592 1051 1604 1085
rect 1638 1051 1650 1085
rect 1592 1017 1650 1051
rect 1592 983 1604 1017
rect 1638 983 1650 1017
rect 1592 949 1650 983
rect 1592 915 1604 949
rect 1638 915 1650 949
rect 1592 881 1650 915
rect 1592 847 1604 881
rect 1638 847 1650 881
rect 1592 813 1650 847
rect 1592 779 1604 813
rect 1638 779 1650 813
rect 1592 745 1650 779
rect 1592 711 1604 745
rect 1638 711 1650 745
rect 1592 677 1650 711
rect 1592 643 1604 677
rect 1638 643 1650 677
rect 1592 600 1650 643
rect 2050 1357 2108 1400
rect 2050 1323 2062 1357
rect 2096 1323 2108 1357
rect 2050 1289 2108 1323
rect 2050 1255 2062 1289
rect 2096 1255 2108 1289
rect 2050 1221 2108 1255
rect 2050 1187 2062 1221
rect 2096 1187 2108 1221
rect 2050 1153 2108 1187
rect 2050 1119 2062 1153
rect 2096 1119 2108 1153
rect 2050 1085 2108 1119
rect 2050 1051 2062 1085
rect 2096 1051 2108 1085
rect 2050 1017 2108 1051
rect 2050 983 2062 1017
rect 2096 983 2108 1017
rect 2050 949 2108 983
rect 2050 915 2062 949
rect 2096 915 2108 949
rect 2050 881 2108 915
rect 2050 847 2062 881
rect 2096 847 2108 881
rect 2050 813 2108 847
rect 2050 779 2062 813
rect 2096 779 2108 813
rect 2050 745 2108 779
rect 2050 711 2062 745
rect 2096 711 2108 745
rect 2050 677 2108 711
rect 2050 643 2062 677
rect 2096 643 2108 677
rect 2050 600 2108 643
rect 2508 1357 2566 1400
rect 2508 1323 2520 1357
rect 2554 1323 2566 1357
rect 2508 1289 2566 1323
rect 2508 1255 2520 1289
rect 2554 1255 2566 1289
rect 2508 1221 2566 1255
rect 2508 1187 2520 1221
rect 2554 1187 2566 1221
rect 2508 1153 2566 1187
rect 2508 1119 2520 1153
rect 2554 1119 2566 1153
rect 2508 1085 2566 1119
rect 2508 1051 2520 1085
rect 2554 1051 2566 1085
rect 2508 1017 2566 1051
rect 2508 983 2520 1017
rect 2554 983 2566 1017
rect 2508 949 2566 983
rect 2508 915 2520 949
rect 2554 915 2566 949
rect 2508 881 2566 915
rect 2508 847 2520 881
rect 2554 847 2566 881
rect 2508 813 2566 847
rect 2508 779 2520 813
rect 2554 779 2566 813
rect 2508 745 2566 779
rect 2508 711 2520 745
rect 2554 711 2566 745
rect 2508 677 2566 711
rect 2508 643 2520 677
rect 2554 643 2566 677
rect 2508 600 2566 643
rect 2966 1357 3024 1400
rect 2966 1323 2978 1357
rect 3012 1323 3024 1357
rect 2966 1289 3024 1323
rect 2966 1255 2978 1289
rect 3012 1255 3024 1289
rect 2966 1221 3024 1255
rect 2966 1187 2978 1221
rect 3012 1187 3024 1221
rect 2966 1153 3024 1187
rect 2966 1119 2978 1153
rect 3012 1119 3024 1153
rect 2966 1085 3024 1119
rect 2966 1051 2978 1085
rect 3012 1051 3024 1085
rect 2966 1017 3024 1051
rect 2966 983 2978 1017
rect 3012 983 3024 1017
rect 2966 949 3024 983
rect 2966 915 2978 949
rect 3012 915 3024 949
rect 2966 881 3024 915
rect 2966 847 2978 881
rect 3012 847 3024 881
rect 2966 813 3024 847
rect 2966 779 2978 813
rect 3012 779 3024 813
rect 2966 745 3024 779
rect 2966 711 2978 745
rect 3012 711 3024 745
rect 2966 677 3024 711
rect 2966 643 2978 677
rect 3012 643 3024 677
rect 2966 600 3024 643
rect 3424 1357 3482 1400
rect 3424 1323 3436 1357
rect 3470 1323 3482 1357
rect 3424 1289 3482 1323
rect 3424 1255 3436 1289
rect 3470 1255 3482 1289
rect 3424 1221 3482 1255
rect 3424 1187 3436 1221
rect 3470 1187 3482 1221
rect 3424 1153 3482 1187
rect 3424 1119 3436 1153
rect 3470 1119 3482 1153
rect 3424 1085 3482 1119
rect 3424 1051 3436 1085
rect 3470 1051 3482 1085
rect 3424 1017 3482 1051
rect 3424 983 3436 1017
rect 3470 983 3482 1017
rect 3424 949 3482 983
rect 3424 915 3436 949
rect 3470 915 3482 949
rect 3424 881 3482 915
rect 3424 847 3436 881
rect 3470 847 3482 881
rect 3424 813 3482 847
rect 3424 779 3436 813
rect 3470 779 3482 813
rect 3424 745 3482 779
rect 3424 711 3436 745
rect 3470 711 3482 745
rect 3424 677 3482 711
rect 3424 643 3436 677
rect 3470 643 3482 677
rect 3424 600 3482 643
rect 3882 1357 3940 1400
rect 3882 1323 3894 1357
rect 3928 1323 3940 1357
rect 3882 1289 3940 1323
rect 3882 1255 3894 1289
rect 3928 1255 3940 1289
rect 3882 1221 3940 1255
rect 3882 1187 3894 1221
rect 3928 1187 3940 1221
rect 3882 1153 3940 1187
rect 3882 1119 3894 1153
rect 3928 1119 3940 1153
rect 3882 1085 3940 1119
rect 3882 1051 3894 1085
rect 3928 1051 3940 1085
rect 3882 1017 3940 1051
rect 3882 983 3894 1017
rect 3928 983 3940 1017
rect 3882 949 3940 983
rect 3882 915 3894 949
rect 3928 915 3940 949
rect 3882 881 3940 915
rect 3882 847 3894 881
rect 3928 847 3940 881
rect 3882 813 3940 847
rect 3882 779 3894 813
rect 3928 779 3940 813
rect 3882 745 3940 779
rect 3882 711 3894 745
rect 3928 711 3940 745
rect 3882 677 3940 711
rect 3882 643 3894 677
rect 3928 643 3940 677
rect 3882 600 3940 643
rect 4340 1357 4398 1400
rect 4340 1323 4352 1357
rect 4386 1323 4398 1357
rect 4340 1289 4398 1323
rect 4340 1255 4352 1289
rect 4386 1255 4398 1289
rect 4340 1221 4398 1255
rect 4340 1187 4352 1221
rect 4386 1187 4398 1221
rect 4340 1153 4398 1187
rect 4340 1119 4352 1153
rect 4386 1119 4398 1153
rect 4340 1085 4398 1119
rect 4340 1051 4352 1085
rect 4386 1051 4398 1085
rect 4340 1017 4398 1051
rect 4340 983 4352 1017
rect 4386 983 4398 1017
rect 4340 949 4398 983
rect 4340 915 4352 949
rect 4386 915 4398 949
rect 4340 881 4398 915
rect 4340 847 4352 881
rect 4386 847 4398 881
rect 4340 813 4398 847
rect 4340 779 4352 813
rect 4386 779 4398 813
rect 4340 745 4398 779
rect 4340 711 4352 745
rect 4386 711 4398 745
rect 4340 677 4398 711
rect 4340 643 4352 677
rect 4386 643 4398 677
rect 4340 600 4398 643
<< ndiffc >>
rect 230 1323 264 1357
rect 230 1255 264 1289
rect 230 1187 264 1221
rect 230 1119 264 1153
rect 230 1051 264 1085
rect 230 983 264 1017
rect 230 915 264 949
rect 230 847 264 881
rect 230 779 264 813
rect 230 711 264 745
rect 230 643 264 677
rect 688 1323 722 1357
rect 688 1255 722 1289
rect 688 1187 722 1221
rect 688 1119 722 1153
rect 688 1051 722 1085
rect 688 983 722 1017
rect 688 915 722 949
rect 688 847 722 881
rect 688 779 722 813
rect 688 711 722 745
rect 688 643 722 677
rect 1146 1323 1180 1357
rect 1146 1255 1180 1289
rect 1146 1187 1180 1221
rect 1146 1119 1180 1153
rect 1146 1051 1180 1085
rect 1146 983 1180 1017
rect 1146 915 1180 949
rect 1146 847 1180 881
rect 1146 779 1180 813
rect 1146 711 1180 745
rect 1146 643 1180 677
rect 1604 1323 1638 1357
rect 1604 1255 1638 1289
rect 1604 1187 1638 1221
rect 1604 1119 1638 1153
rect 1604 1051 1638 1085
rect 1604 983 1638 1017
rect 1604 915 1638 949
rect 1604 847 1638 881
rect 1604 779 1638 813
rect 1604 711 1638 745
rect 1604 643 1638 677
rect 2062 1323 2096 1357
rect 2062 1255 2096 1289
rect 2062 1187 2096 1221
rect 2062 1119 2096 1153
rect 2062 1051 2096 1085
rect 2062 983 2096 1017
rect 2062 915 2096 949
rect 2062 847 2096 881
rect 2062 779 2096 813
rect 2062 711 2096 745
rect 2062 643 2096 677
rect 2520 1323 2554 1357
rect 2520 1255 2554 1289
rect 2520 1187 2554 1221
rect 2520 1119 2554 1153
rect 2520 1051 2554 1085
rect 2520 983 2554 1017
rect 2520 915 2554 949
rect 2520 847 2554 881
rect 2520 779 2554 813
rect 2520 711 2554 745
rect 2520 643 2554 677
rect 2978 1323 3012 1357
rect 2978 1255 3012 1289
rect 2978 1187 3012 1221
rect 2978 1119 3012 1153
rect 2978 1051 3012 1085
rect 2978 983 3012 1017
rect 2978 915 3012 949
rect 2978 847 3012 881
rect 2978 779 3012 813
rect 2978 711 3012 745
rect 2978 643 3012 677
rect 3436 1323 3470 1357
rect 3436 1255 3470 1289
rect 3436 1187 3470 1221
rect 3436 1119 3470 1153
rect 3436 1051 3470 1085
rect 3436 983 3470 1017
rect 3436 915 3470 949
rect 3436 847 3470 881
rect 3436 779 3470 813
rect 3436 711 3470 745
rect 3436 643 3470 677
rect 3894 1323 3928 1357
rect 3894 1255 3928 1289
rect 3894 1187 3928 1221
rect 3894 1119 3928 1153
rect 3894 1051 3928 1085
rect 3894 983 3928 1017
rect 3894 915 3928 949
rect 3894 847 3928 881
rect 3894 779 3928 813
rect 3894 711 3928 745
rect 3894 643 3928 677
rect 4352 1323 4386 1357
rect 4352 1255 4386 1289
rect 4352 1187 4386 1221
rect 4352 1119 4386 1153
rect 4352 1051 4386 1085
rect 4352 983 4386 1017
rect 4352 915 4386 949
rect 4352 847 4386 881
rect 4352 779 4386 813
rect 4352 711 4386 745
rect 4352 643 4386 677
<< psubdiff >>
rect 158 157 198 200
rect 158 123 161 157
rect 195 123 198 157
rect 158 80 198 123
rect 1218 127 1338 130
rect 1218 93 1263 127
rect 1297 93 1338 127
rect 1218 80 1338 93
rect 2518 127 2638 130
rect 2518 93 2563 127
rect 2597 93 2638 127
rect 2518 80 2638 93
<< psubdiffcont >>
rect 161 123 195 157
rect 1263 93 1297 127
rect 2563 93 2597 127
<< poly >>
rect 276 1400 676 1426
rect 734 1400 1134 1426
rect 1192 1400 1592 1426
rect 1650 1400 2050 1426
rect 2108 1400 2508 1426
rect 2566 1400 2966 1426
rect 3024 1400 3424 1426
rect 3482 1400 3882 1426
rect 3940 1400 4340 1426
rect 276 574 676 600
rect 734 574 1134 600
rect 1192 574 1592 600
rect 1650 574 2050 600
rect 2108 574 2508 600
rect 2566 574 2966 600
rect 3024 574 3424 600
rect 3482 574 3882 600
rect 3940 574 4340 600
rect 424 384 544 574
rect 880 384 1000 574
rect 1336 384 1456 574
rect 1792 384 1912 574
rect 2248 384 2368 574
rect 2704 384 2824 574
rect 3160 384 3280 574
rect 3616 384 3736 574
rect 4072 384 4192 574
rect 298 351 4398 384
rect 298 317 401 351
rect 435 317 801 351
rect 835 317 1201 351
rect 1235 317 1601 351
rect 1635 317 2001 351
rect 2035 317 2401 351
rect 2435 317 2801 351
rect 2835 317 3201 351
rect 3235 317 3601 351
rect 3635 317 4001 351
rect 4035 317 4398 351
rect 298 284 4398 317
<< polycont >>
rect 401 317 435 351
rect 801 317 835 351
rect 1201 317 1235 351
rect 1601 317 1635 351
rect 2001 317 2035 351
rect 2401 317 2435 351
rect 2801 317 2835 351
rect 3201 317 3235 351
rect 3601 317 3635 351
rect 4001 317 4035 351
<< locali >>
rect 120 1897 4398 1910
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3201 1897
rect 3235 1863 3601 1897
rect 3635 1863 4001 1897
rect 4035 1863 4398 1897
rect 120 1850 4398 1863
rect 218 1690 4398 1750
rect 687 1404 721 1690
rect 1603 1404 1637 1690
rect 2519 1404 2553 1690
rect 3435 1404 3469 1690
rect 4351 1404 4385 1690
rect 230 1377 264 1404
rect 687 1386 722 1404
rect 230 1305 264 1323
rect 230 1233 264 1255
rect 230 1161 264 1187
rect 230 1089 264 1119
rect 230 1017 264 1051
rect 230 949 264 983
rect 230 881 264 911
rect 230 813 264 839
rect 230 745 264 767
rect 230 677 264 695
rect 229 623 230 654
rect 229 596 264 623
rect 688 1377 722 1386
rect 688 1305 722 1323
rect 688 1233 722 1255
rect 688 1161 722 1187
rect 688 1089 722 1119
rect 688 1017 722 1051
rect 688 949 722 983
rect 688 881 722 911
rect 688 813 722 839
rect 688 745 722 767
rect 688 677 722 695
rect 1146 1377 1180 1404
rect 1603 1386 1638 1404
rect 1146 1305 1180 1323
rect 1146 1233 1180 1255
rect 1146 1161 1180 1187
rect 1146 1089 1180 1119
rect 1146 1017 1180 1051
rect 1146 949 1180 983
rect 1146 881 1180 911
rect 1146 813 1180 839
rect 1146 745 1180 767
rect 1146 677 1180 695
rect 688 596 722 623
rect 1145 623 1146 654
rect 1145 596 1180 623
rect 1604 1377 1638 1386
rect 1604 1305 1638 1323
rect 1604 1233 1638 1255
rect 1604 1161 1638 1187
rect 1604 1089 1638 1119
rect 1604 1017 1638 1051
rect 1604 949 1638 983
rect 1604 881 1638 911
rect 1604 813 1638 839
rect 1604 745 1638 767
rect 1604 677 1638 695
rect 2062 1377 2096 1404
rect 2519 1386 2554 1404
rect 2062 1305 2096 1323
rect 2062 1233 2096 1255
rect 2062 1161 2096 1187
rect 2062 1089 2096 1119
rect 2062 1017 2096 1051
rect 2062 949 2096 983
rect 2062 881 2096 911
rect 2062 813 2096 839
rect 2062 745 2096 767
rect 2062 677 2096 695
rect 1604 596 1638 623
rect 2061 623 2062 654
rect 2061 596 2096 623
rect 2520 1377 2554 1386
rect 2520 1305 2554 1323
rect 2520 1233 2554 1255
rect 2520 1161 2554 1187
rect 2520 1089 2554 1119
rect 2520 1017 2554 1051
rect 2520 949 2554 983
rect 2520 881 2554 911
rect 2520 813 2554 839
rect 2520 745 2554 767
rect 2520 677 2554 695
rect 2978 1377 3012 1404
rect 3435 1386 3470 1404
rect 2978 1305 3012 1323
rect 2978 1233 3012 1255
rect 2978 1161 3012 1187
rect 2978 1089 3012 1119
rect 2978 1017 3012 1051
rect 2978 949 3012 983
rect 2978 881 3012 911
rect 2978 813 3012 839
rect 2978 745 3012 767
rect 2978 677 3012 695
rect 2520 596 2554 623
rect 2977 623 2978 654
rect 2977 596 3012 623
rect 3436 1377 3470 1386
rect 3436 1305 3470 1323
rect 3436 1233 3470 1255
rect 3436 1161 3470 1187
rect 3436 1089 3470 1119
rect 3436 1017 3470 1051
rect 3436 949 3470 983
rect 3436 881 3470 911
rect 3436 813 3470 839
rect 3436 745 3470 767
rect 3436 677 3470 695
rect 3894 1377 3928 1404
rect 4351 1386 4386 1404
rect 3894 1305 3928 1323
rect 3894 1233 3928 1255
rect 3894 1161 3928 1187
rect 3894 1089 3928 1119
rect 3894 1017 3928 1051
rect 3894 949 3928 983
rect 3894 881 3928 911
rect 3894 813 3928 839
rect 3894 745 3928 767
rect 3894 677 3928 695
rect 3436 596 3470 623
rect 3893 623 3894 654
rect 3893 596 3928 623
rect 4352 1377 4386 1386
rect 4352 1305 4386 1323
rect 4352 1233 4386 1255
rect 4352 1161 4386 1187
rect 4352 1089 4386 1119
rect 4352 1017 4386 1051
rect 4352 949 4386 983
rect 4352 881 4386 911
rect 4352 813 4386 839
rect 4352 745 4386 767
rect 4352 677 4386 695
rect 4352 596 4386 623
rect 229 530 263 596
rect 1145 530 1179 596
rect 2061 530 2095 596
rect 2977 530 3011 596
rect 3893 530 3927 596
rect 218 470 4398 530
rect 298 351 4398 364
rect 298 317 401 351
rect 435 317 801 351
rect 835 317 1201 351
rect 1235 317 1601 351
rect 1635 317 2001 351
rect 2035 317 2401 351
rect 2435 317 2801 351
rect 2835 317 3201 351
rect 3235 317 3601 351
rect 3635 317 4001 351
rect 4035 317 4398 351
rect 298 304 4398 317
rect 148 157 208 240
rect 148 123 161 157
rect 195 123 208 157
rect 148 30 208 123
rect 1198 127 1358 150
rect 1198 93 1263 127
rect 1297 93 1358 127
rect 1198 30 1358 93
rect 2498 127 2658 150
rect 2498 93 2563 127
rect 2597 93 2658 127
rect 2498 30 2658 93
rect 120 17 4398 30
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3201 17
rect 3235 -17 3601 17
rect 3635 -17 4001 17
rect 4035 -17 4398 17
rect 120 -30 4398 -17
<< viali >>
rect 401 1863 435 1897
rect 801 1863 835 1897
rect 1201 1863 1235 1897
rect 1601 1863 1635 1897
rect 2001 1863 2035 1897
rect 2401 1863 2435 1897
rect 2801 1863 2835 1897
rect 3201 1863 3235 1897
rect 3601 1863 3635 1897
rect 4001 1863 4035 1897
rect 230 1357 264 1377
rect 230 1343 264 1357
rect 230 1289 264 1305
rect 230 1271 264 1289
rect 230 1221 264 1233
rect 230 1199 264 1221
rect 230 1153 264 1161
rect 230 1127 264 1153
rect 230 1085 264 1089
rect 230 1055 264 1085
rect 230 983 264 1017
rect 230 915 264 945
rect 230 911 264 915
rect 230 847 264 873
rect 230 839 264 847
rect 230 779 264 801
rect 230 767 264 779
rect 230 711 264 729
rect 230 695 264 711
rect 230 643 264 657
rect 230 623 264 643
rect 688 1357 722 1377
rect 688 1343 722 1357
rect 688 1289 722 1305
rect 688 1271 722 1289
rect 688 1221 722 1233
rect 688 1199 722 1221
rect 688 1153 722 1161
rect 688 1127 722 1153
rect 688 1085 722 1089
rect 688 1055 722 1085
rect 688 983 722 1017
rect 688 915 722 945
rect 688 911 722 915
rect 688 847 722 873
rect 688 839 722 847
rect 688 779 722 801
rect 688 767 722 779
rect 688 711 722 729
rect 688 695 722 711
rect 688 643 722 657
rect 1146 1357 1180 1377
rect 1146 1343 1180 1357
rect 1146 1289 1180 1305
rect 1146 1271 1180 1289
rect 1146 1221 1180 1233
rect 1146 1199 1180 1221
rect 1146 1153 1180 1161
rect 1146 1127 1180 1153
rect 1146 1085 1180 1089
rect 1146 1055 1180 1085
rect 1146 983 1180 1017
rect 1146 915 1180 945
rect 1146 911 1180 915
rect 1146 847 1180 873
rect 1146 839 1180 847
rect 1146 779 1180 801
rect 1146 767 1180 779
rect 1146 711 1180 729
rect 1146 695 1180 711
rect 688 623 722 643
rect 1146 643 1180 657
rect 1146 623 1180 643
rect 1604 1357 1638 1377
rect 1604 1343 1638 1357
rect 1604 1289 1638 1305
rect 1604 1271 1638 1289
rect 1604 1221 1638 1233
rect 1604 1199 1638 1221
rect 1604 1153 1638 1161
rect 1604 1127 1638 1153
rect 1604 1085 1638 1089
rect 1604 1055 1638 1085
rect 1604 983 1638 1017
rect 1604 915 1638 945
rect 1604 911 1638 915
rect 1604 847 1638 873
rect 1604 839 1638 847
rect 1604 779 1638 801
rect 1604 767 1638 779
rect 1604 711 1638 729
rect 1604 695 1638 711
rect 1604 643 1638 657
rect 2062 1357 2096 1377
rect 2062 1343 2096 1357
rect 2062 1289 2096 1305
rect 2062 1271 2096 1289
rect 2062 1221 2096 1233
rect 2062 1199 2096 1221
rect 2062 1153 2096 1161
rect 2062 1127 2096 1153
rect 2062 1085 2096 1089
rect 2062 1055 2096 1085
rect 2062 983 2096 1017
rect 2062 915 2096 945
rect 2062 911 2096 915
rect 2062 847 2096 873
rect 2062 839 2096 847
rect 2062 779 2096 801
rect 2062 767 2096 779
rect 2062 711 2096 729
rect 2062 695 2096 711
rect 1604 623 1638 643
rect 2062 643 2096 657
rect 2062 623 2096 643
rect 2520 1357 2554 1377
rect 2520 1343 2554 1357
rect 2520 1289 2554 1305
rect 2520 1271 2554 1289
rect 2520 1221 2554 1233
rect 2520 1199 2554 1221
rect 2520 1153 2554 1161
rect 2520 1127 2554 1153
rect 2520 1085 2554 1089
rect 2520 1055 2554 1085
rect 2520 983 2554 1017
rect 2520 915 2554 945
rect 2520 911 2554 915
rect 2520 847 2554 873
rect 2520 839 2554 847
rect 2520 779 2554 801
rect 2520 767 2554 779
rect 2520 711 2554 729
rect 2520 695 2554 711
rect 2520 643 2554 657
rect 2978 1357 3012 1377
rect 2978 1343 3012 1357
rect 2978 1289 3012 1305
rect 2978 1271 3012 1289
rect 2978 1221 3012 1233
rect 2978 1199 3012 1221
rect 2978 1153 3012 1161
rect 2978 1127 3012 1153
rect 2978 1085 3012 1089
rect 2978 1055 3012 1085
rect 2978 983 3012 1017
rect 2978 915 3012 945
rect 2978 911 3012 915
rect 2978 847 3012 873
rect 2978 839 3012 847
rect 2978 779 3012 801
rect 2978 767 3012 779
rect 2978 711 3012 729
rect 2978 695 3012 711
rect 2520 623 2554 643
rect 2978 643 3012 657
rect 2978 623 3012 643
rect 3436 1357 3470 1377
rect 3436 1343 3470 1357
rect 3436 1289 3470 1305
rect 3436 1271 3470 1289
rect 3436 1221 3470 1233
rect 3436 1199 3470 1221
rect 3436 1153 3470 1161
rect 3436 1127 3470 1153
rect 3436 1085 3470 1089
rect 3436 1055 3470 1085
rect 3436 983 3470 1017
rect 3436 915 3470 945
rect 3436 911 3470 915
rect 3436 847 3470 873
rect 3436 839 3470 847
rect 3436 779 3470 801
rect 3436 767 3470 779
rect 3436 711 3470 729
rect 3436 695 3470 711
rect 3436 643 3470 657
rect 3894 1357 3928 1377
rect 3894 1343 3928 1357
rect 3894 1289 3928 1305
rect 3894 1271 3928 1289
rect 3894 1221 3928 1233
rect 3894 1199 3928 1221
rect 3894 1153 3928 1161
rect 3894 1127 3928 1153
rect 3894 1085 3928 1089
rect 3894 1055 3928 1085
rect 3894 983 3928 1017
rect 3894 915 3928 945
rect 3894 911 3928 915
rect 3894 847 3928 873
rect 3894 839 3928 847
rect 3894 779 3928 801
rect 3894 767 3928 779
rect 3894 711 3928 729
rect 3894 695 3928 711
rect 3436 623 3470 643
rect 3894 643 3928 657
rect 3894 623 3928 643
rect 4352 1357 4386 1377
rect 4352 1343 4386 1357
rect 4352 1289 4386 1305
rect 4352 1271 4386 1289
rect 4352 1221 4386 1233
rect 4352 1199 4386 1221
rect 4352 1153 4386 1161
rect 4352 1127 4386 1153
rect 4352 1085 4386 1089
rect 4352 1055 4386 1085
rect 4352 983 4386 1017
rect 4352 915 4386 945
rect 4352 911 4386 915
rect 4352 847 4386 873
rect 4352 839 4386 847
rect 4352 779 4386 801
rect 4352 767 4386 779
rect 4352 711 4386 729
rect 4352 695 4386 711
rect 4352 643 4386 657
rect 4352 623 4386 643
rect 401 -17 435 17
rect 801 -17 835 17
rect 1201 -17 1235 17
rect 1601 -17 1635 17
rect 2001 -17 2035 17
rect 2401 -17 2435 17
rect 2801 -17 2835 17
rect 3201 -17 3235 17
rect 3601 -17 3635 17
rect 4001 -17 4035 17
<< metal1 >>
rect 120 1897 4398 1940
rect 120 1863 401 1897
rect 435 1863 801 1897
rect 835 1863 1201 1897
rect 1235 1863 1601 1897
rect 1635 1863 2001 1897
rect 2035 1863 2401 1897
rect 2435 1863 2801 1897
rect 2835 1863 3201 1897
rect 3235 1863 3601 1897
rect 3635 1863 4001 1897
rect 4035 1863 4398 1897
rect 120 1820 4398 1863
rect 224 1377 270 1400
rect 224 1343 230 1377
rect 264 1343 270 1377
rect 224 1305 270 1343
rect 224 1271 230 1305
rect 264 1271 270 1305
rect 224 1233 270 1271
rect 224 1199 230 1233
rect 264 1199 270 1233
rect 224 1161 270 1199
rect 224 1127 230 1161
rect 264 1127 270 1161
rect 224 1089 270 1127
rect 224 1055 230 1089
rect 264 1055 270 1089
rect 224 1017 270 1055
rect 224 983 230 1017
rect 264 983 270 1017
rect 224 945 270 983
rect 224 911 230 945
rect 264 911 270 945
rect 224 873 270 911
rect 224 839 230 873
rect 264 839 270 873
rect 224 801 270 839
rect 224 767 230 801
rect 264 767 270 801
rect 224 729 270 767
rect 224 695 230 729
rect 264 695 270 729
rect 224 657 270 695
rect 224 623 230 657
rect 264 623 270 657
rect 224 600 270 623
rect 682 1377 728 1400
rect 682 1343 688 1377
rect 722 1343 728 1377
rect 682 1305 728 1343
rect 682 1271 688 1305
rect 722 1271 728 1305
rect 682 1233 728 1271
rect 682 1199 688 1233
rect 722 1199 728 1233
rect 682 1161 728 1199
rect 682 1127 688 1161
rect 722 1127 728 1161
rect 682 1089 728 1127
rect 682 1055 688 1089
rect 722 1055 728 1089
rect 682 1017 728 1055
rect 682 983 688 1017
rect 722 983 728 1017
rect 682 945 728 983
rect 682 911 688 945
rect 722 911 728 945
rect 682 873 728 911
rect 682 839 688 873
rect 722 839 728 873
rect 682 801 728 839
rect 682 767 688 801
rect 722 767 728 801
rect 682 729 728 767
rect 682 695 688 729
rect 722 695 728 729
rect 682 657 728 695
rect 682 623 688 657
rect 722 623 728 657
rect 682 600 728 623
rect 1140 1377 1186 1400
rect 1140 1343 1146 1377
rect 1180 1343 1186 1377
rect 1140 1305 1186 1343
rect 1140 1271 1146 1305
rect 1180 1271 1186 1305
rect 1140 1233 1186 1271
rect 1140 1199 1146 1233
rect 1180 1199 1186 1233
rect 1140 1161 1186 1199
rect 1140 1127 1146 1161
rect 1180 1127 1186 1161
rect 1140 1089 1186 1127
rect 1140 1055 1146 1089
rect 1180 1055 1186 1089
rect 1140 1017 1186 1055
rect 1140 983 1146 1017
rect 1180 983 1186 1017
rect 1140 945 1186 983
rect 1140 911 1146 945
rect 1180 911 1186 945
rect 1140 873 1186 911
rect 1140 839 1146 873
rect 1180 839 1186 873
rect 1140 801 1186 839
rect 1140 767 1146 801
rect 1180 767 1186 801
rect 1140 729 1186 767
rect 1140 695 1146 729
rect 1180 695 1186 729
rect 1140 657 1186 695
rect 1140 623 1146 657
rect 1180 623 1186 657
rect 1140 600 1186 623
rect 1598 1377 1644 1400
rect 1598 1343 1604 1377
rect 1638 1343 1644 1377
rect 1598 1305 1644 1343
rect 1598 1271 1604 1305
rect 1638 1271 1644 1305
rect 1598 1233 1644 1271
rect 1598 1199 1604 1233
rect 1638 1199 1644 1233
rect 1598 1161 1644 1199
rect 1598 1127 1604 1161
rect 1638 1127 1644 1161
rect 1598 1089 1644 1127
rect 1598 1055 1604 1089
rect 1638 1055 1644 1089
rect 1598 1017 1644 1055
rect 1598 983 1604 1017
rect 1638 983 1644 1017
rect 1598 945 1644 983
rect 1598 911 1604 945
rect 1638 911 1644 945
rect 1598 873 1644 911
rect 1598 839 1604 873
rect 1638 839 1644 873
rect 1598 801 1644 839
rect 1598 767 1604 801
rect 1638 767 1644 801
rect 1598 729 1644 767
rect 1598 695 1604 729
rect 1638 695 1644 729
rect 1598 657 1644 695
rect 1598 623 1604 657
rect 1638 623 1644 657
rect 1598 600 1644 623
rect 2056 1377 2102 1400
rect 2056 1343 2062 1377
rect 2096 1343 2102 1377
rect 2056 1305 2102 1343
rect 2056 1271 2062 1305
rect 2096 1271 2102 1305
rect 2056 1233 2102 1271
rect 2056 1199 2062 1233
rect 2096 1199 2102 1233
rect 2056 1161 2102 1199
rect 2056 1127 2062 1161
rect 2096 1127 2102 1161
rect 2056 1089 2102 1127
rect 2056 1055 2062 1089
rect 2096 1055 2102 1089
rect 2056 1017 2102 1055
rect 2056 983 2062 1017
rect 2096 983 2102 1017
rect 2056 945 2102 983
rect 2056 911 2062 945
rect 2096 911 2102 945
rect 2056 873 2102 911
rect 2056 839 2062 873
rect 2096 839 2102 873
rect 2056 801 2102 839
rect 2056 767 2062 801
rect 2096 767 2102 801
rect 2056 729 2102 767
rect 2056 695 2062 729
rect 2096 695 2102 729
rect 2056 657 2102 695
rect 2056 623 2062 657
rect 2096 623 2102 657
rect 2056 600 2102 623
rect 2514 1377 2560 1400
rect 2514 1343 2520 1377
rect 2554 1343 2560 1377
rect 2514 1305 2560 1343
rect 2514 1271 2520 1305
rect 2554 1271 2560 1305
rect 2514 1233 2560 1271
rect 2514 1199 2520 1233
rect 2554 1199 2560 1233
rect 2514 1161 2560 1199
rect 2514 1127 2520 1161
rect 2554 1127 2560 1161
rect 2514 1089 2560 1127
rect 2514 1055 2520 1089
rect 2554 1055 2560 1089
rect 2514 1017 2560 1055
rect 2514 983 2520 1017
rect 2554 983 2560 1017
rect 2514 945 2560 983
rect 2514 911 2520 945
rect 2554 911 2560 945
rect 2514 873 2560 911
rect 2514 839 2520 873
rect 2554 839 2560 873
rect 2514 801 2560 839
rect 2514 767 2520 801
rect 2554 767 2560 801
rect 2514 729 2560 767
rect 2514 695 2520 729
rect 2554 695 2560 729
rect 2514 657 2560 695
rect 2514 623 2520 657
rect 2554 623 2560 657
rect 2514 600 2560 623
rect 2972 1377 3018 1400
rect 2972 1343 2978 1377
rect 3012 1343 3018 1377
rect 2972 1305 3018 1343
rect 2972 1271 2978 1305
rect 3012 1271 3018 1305
rect 2972 1233 3018 1271
rect 2972 1199 2978 1233
rect 3012 1199 3018 1233
rect 2972 1161 3018 1199
rect 2972 1127 2978 1161
rect 3012 1127 3018 1161
rect 2972 1089 3018 1127
rect 2972 1055 2978 1089
rect 3012 1055 3018 1089
rect 2972 1017 3018 1055
rect 2972 983 2978 1017
rect 3012 983 3018 1017
rect 2972 945 3018 983
rect 2972 911 2978 945
rect 3012 911 3018 945
rect 2972 873 3018 911
rect 2972 839 2978 873
rect 3012 839 3018 873
rect 2972 801 3018 839
rect 2972 767 2978 801
rect 3012 767 3018 801
rect 2972 729 3018 767
rect 2972 695 2978 729
rect 3012 695 3018 729
rect 2972 657 3018 695
rect 2972 623 2978 657
rect 3012 623 3018 657
rect 2972 600 3018 623
rect 3430 1377 3476 1400
rect 3430 1343 3436 1377
rect 3470 1343 3476 1377
rect 3430 1305 3476 1343
rect 3430 1271 3436 1305
rect 3470 1271 3476 1305
rect 3430 1233 3476 1271
rect 3430 1199 3436 1233
rect 3470 1199 3476 1233
rect 3430 1161 3476 1199
rect 3430 1127 3436 1161
rect 3470 1127 3476 1161
rect 3430 1089 3476 1127
rect 3430 1055 3436 1089
rect 3470 1055 3476 1089
rect 3430 1017 3476 1055
rect 3430 983 3436 1017
rect 3470 983 3476 1017
rect 3430 945 3476 983
rect 3430 911 3436 945
rect 3470 911 3476 945
rect 3430 873 3476 911
rect 3430 839 3436 873
rect 3470 839 3476 873
rect 3430 801 3476 839
rect 3430 767 3436 801
rect 3470 767 3476 801
rect 3430 729 3476 767
rect 3430 695 3436 729
rect 3470 695 3476 729
rect 3430 657 3476 695
rect 3430 623 3436 657
rect 3470 623 3476 657
rect 3430 600 3476 623
rect 3888 1377 3934 1400
rect 3888 1343 3894 1377
rect 3928 1343 3934 1377
rect 3888 1305 3934 1343
rect 3888 1271 3894 1305
rect 3928 1271 3934 1305
rect 3888 1233 3934 1271
rect 3888 1199 3894 1233
rect 3928 1199 3934 1233
rect 3888 1161 3934 1199
rect 3888 1127 3894 1161
rect 3928 1127 3934 1161
rect 3888 1089 3934 1127
rect 3888 1055 3894 1089
rect 3928 1055 3934 1089
rect 3888 1017 3934 1055
rect 3888 983 3894 1017
rect 3928 983 3934 1017
rect 3888 945 3934 983
rect 3888 911 3894 945
rect 3928 911 3934 945
rect 3888 873 3934 911
rect 3888 839 3894 873
rect 3928 839 3934 873
rect 3888 801 3934 839
rect 3888 767 3894 801
rect 3928 767 3934 801
rect 3888 729 3934 767
rect 3888 695 3894 729
rect 3928 695 3934 729
rect 3888 657 3934 695
rect 3888 623 3894 657
rect 3928 623 3934 657
rect 3888 600 3934 623
rect 4346 1377 4392 1400
rect 4346 1343 4352 1377
rect 4386 1343 4392 1377
rect 4346 1305 4392 1343
rect 4346 1271 4352 1305
rect 4386 1271 4392 1305
rect 4346 1233 4392 1271
rect 4346 1199 4352 1233
rect 4386 1199 4392 1233
rect 4346 1161 4392 1199
rect 4346 1127 4352 1161
rect 4386 1127 4392 1161
rect 4346 1089 4392 1127
rect 4346 1055 4352 1089
rect 4386 1055 4392 1089
rect 4346 1017 4392 1055
rect 4346 983 4352 1017
rect 4386 983 4392 1017
rect 4346 945 4392 983
rect 4346 911 4352 945
rect 4386 911 4392 945
rect 4346 873 4392 911
rect 4346 839 4352 873
rect 4386 839 4392 873
rect 4346 801 4392 839
rect 4346 767 4352 801
rect 4386 767 4392 801
rect 4346 729 4392 767
rect 4346 695 4352 729
rect 4386 695 4392 729
rect 4346 657 4392 695
rect 4346 623 4352 657
rect 4386 623 4392 657
rect 4346 600 4392 623
rect 120 17 4398 60
rect 120 -17 401 17
rect 435 -17 801 17
rect 835 -17 1201 17
rect 1235 -17 1601 17
rect 1635 -17 2001 17
rect 2035 -17 2401 17
rect 2435 -17 2801 17
rect 2835 -17 3201 17
rect 3235 -17 3601 17
rect 3635 -17 4001 17
rect 4035 -17 4398 17
rect 120 -60 4398 -17
<< labels >>
flabel locali s 4338 304 4398 364 1 FreeSans 1562 0 0 0 GATE
port 1 nsew
flabel locali s 4338 1690 4398 1750 1 FreeSans 1562 0 0 0 SOURCE
port 2 nsew
flabel locali s 4338 470 4398 530 1 FreeSans 1562 0 0 0 DRAIN
port 3 nsew
flabel metal1 s 218 1850 278 1910 1 FreeSans 1562 0 0 0 VPWR
port 4 nsew
flabel metal1 s 218 -30 278 30 1 FreeSans 1562 0 0 0 VGND
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 4518 1880
<< end >>
