magic
tech sky130A
timestamp 1655811994
use bgr_top  bgr_top_0
timestamp 1483682050
transform 1 0 5073 0 1 2958
box 0 0 27278 26418
<< end >>
