magic
tech sky130A
timestamp 1655503347
<< metal2 >>
rect -408 14 408 30
rect -408 -14 -394 14
rect -366 -14 -354 14
rect -326 -14 -314 14
rect -286 -14 -274 14
rect -246 -14 -234 14
rect -206 -14 -194 14
rect -166 -14 -154 14
rect -126 -14 -114 14
rect -86 -14 -74 14
rect -46 -14 -34 14
rect -6 -14 6 14
rect 34 -14 46 14
rect 74 -14 86 14
rect 114 -14 126 14
rect 154 -14 166 14
rect 194 -14 206 14
rect 234 -14 246 14
rect 274 -14 286 14
rect 314 -14 326 14
rect 354 -14 366 14
rect 394 -14 408 14
rect -408 -30 408 -14
<< via2 >>
rect -394 -14 -366 14
rect -354 -14 -326 14
rect -314 -14 -286 14
rect -274 -14 -246 14
rect -234 -14 -206 14
rect -194 -14 -166 14
rect -154 -14 -126 14
rect -114 -14 -86 14
rect -74 -14 -46 14
rect -34 -14 -6 14
rect 6 -14 34 14
rect 46 -14 74 14
rect 86 -14 114 14
rect 126 -14 154 14
rect 166 -14 194 14
rect 206 -14 234 14
rect 246 -14 274 14
rect 286 -14 314 14
rect 326 -14 354 14
rect 366 -14 394 14
<< metal3 >>
rect -408 14 408 30
rect -408 -14 -394 14
rect -366 -14 -354 14
rect -326 -14 -314 14
rect -286 -14 -274 14
rect -246 -14 -234 14
rect -206 -14 -194 14
rect -166 -14 -154 14
rect -126 -14 -114 14
rect -86 -14 -74 14
rect -46 -14 -34 14
rect -6 -14 6 14
rect 34 -14 46 14
rect 74 -14 86 14
rect 114 -14 126 14
rect 154 -14 166 14
rect 194 -14 206 14
rect 234 -14 246 14
rect 274 -14 286 14
rect 314 -14 326 14
rect 354 -14 366 14
rect 394 -14 408 14
rect -408 -30 408 -14
<< end >>
