magic
tech sky130A
magscale 1 2
timestamp 1654901230
<< pwell >>
rect 162 574 730 1426
rect 102 54 194 226
<< nmoslvt >>
rect 246 600 646 1400
<< ndiff >>
rect 188 1357 246 1400
rect 188 1323 200 1357
rect 234 1323 246 1357
rect 188 1289 246 1323
rect 188 1255 200 1289
rect 234 1255 246 1289
rect 188 1221 246 1255
rect 188 1187 200 1221
rect 234 1187 246 1221
rect 188 1153 246 1187
rect 188 1119 200 1153
rect 234 1119 246 1153
rect 188 1085 246 1119
rect 188 1051 200 1085
rect 234 1051 246 1085
rect 188 1017 246 1051
rect 188 983 200 1017
rect 234 983 246 1017
rect 188 949 246 983
rect 188 915 200 949
rect 234 915 246 949
rect 188 881 246 915
rect 188 847 200 881
rect 234 847 246 881
rect 188 813 246 847
rect 188 779 200 813
rect 234 779 246 813
rect 188 745 246 779
rect 188 711 200 745
rect 234 711 246 745
rect 188 677 246 711
rect 188 643 200 677
rect 234 643 246 677
rect 188 600 246 643
rect 646 1357 704 1400
rect 646 1323 658 1357
rect 692 1323 704 1357
rect 646 1289 704 1323
rect 646 1255 658 1289
rect 692 1255 704 1289
rect 646 1221 704 1255
rect 646 1187 658 1221
rect 692 1187 704 1221
rect 646 1153 704 1187
rect 646 1119 658 1153
rect 692 1119 704 1153
rect 646 1085 704 1119
rect 646 1051 658 1085
rect 692 1051 704 1085
rect 646 1017 704 1051
rect 646 983 658 1017
rect 692 983 704 1017
rect 646 949 704 983
rect 646 915 658 949
rect 692 915 704 949
rect 646 881 704 915
rect 646 847 658 881
rect 692 847 704 881
rect 646 813 704 847
rect 646 779 658 813
rect 692 779 704 813
rect 646 745 704 779
rect 646 711 658 745
rect 692 711 704 745
rect 646 677 704 711
rect 646 643 658 677
rect 692 643 704 677
rect 646 600 704 643
<< ndiffc >>
rect 200 1323 234 1357
rect 200 1255 234 1289
rect 200 1187 234 1221
rect 200 1119 234 1153
rect 200 1051 234 1085
rect 200 983 234 1017
rect 200 915 234 949
rect 200 847 234 881
rect 200 779 234 813
rect 200 711 234 745
rect 200 643 234 677
rect 658 1323 692 1357
rect 658 1255 692 1289
rect 658 1187 692 1221
rect 658 1119 692 1153
rect 658 1051 692 1085
rect 658 983 692 1017
rect 658 915 692 949
rect 658 847 692 881
rect 658 779 692 813
rect 658 711 692 745
rect 658 643 692 677
<< psubdiff >>
rect 128 157 168 200
rect 128 123 131 157
rect 165 123 168 157
rect 128 80 168 123
<< psubdiffcont >>
rect 131 123 165 157
<< poly >>
rect 246 1400 646 1426
rect 246 574 646 600
rect 394 224 514 574
rect 268 191 704 224
rect 268 157 371 191
rect 405 157 704 191
rect 268 124 704 157
<< polycont >>
rect 371 157 405 191
<< locali >>
rect 90 1897 704 1910
rect 90 1863 371 1897
rect 405 1863 704 1897
rect 90 1850 704 1863
rect 188 1690 704 1750
rect 657 1404 691 1690
rect 200 1377 234 1404
rect 657 1386 692 1404
rect 200 1305 234 1323
rect 200 1233 234 1255
rect 200 1161 234 1187
rect 200 1089 234 1119
rect 200 1017 234 1051
rect 200 949 234 983
rect 200 881 234 911
rect 200 813 234 839
rect 200 745 234 767
rect 200 677 234 695
rect 199 623 200 654
rect 199 596 234 623
rect 658 1377 692 1386
rect 658 1305 692 1323
rect 658 1233 692 1255
rect 658 1161 692 1187
rect 658 1089 692 1119
rect 658 1017 692 1051
rect 658 949 692 983
rect 658 881 692 911
rect 658 813 692 839
rect 658 745 692 767
rect 658 677 692 695
rect 658 596 692 623
rect 199 430 233 596
rect 188 370 704 430
rect 118 157 178 240
rect 118 123 131 157
rect 165 123 178 157
rect 268 191 704 204
rect 268 157 371 191
rect 405 157 704 191
rect 268 144 704 157
rect 118 30 178 123
rect 90 17 704 30
rect 90 -17 371 17
rect 405 -17 704 17
rect 90 -30 704 -17
<< viali >>
rect 371 1863 405 1897
rect 200 1357 234 1377
rect 200 1343 234 1357
rect 200 1289 234 1305
rect 200 1271 234 1289
rect 200 1221 234 1233
rect 200 1199 234 1221
rect 200 1153 234 1161
rect 200 1127 234 1153
rect 200 1085 234 1089
rect 200 1055 234 1085
rect 200 983 234 1017
rect 200 915 234 945
rect 200 911 234 915
rect 200 847 234 873
rect 200 839 234 847
rect 200 779 234 801
rect 200 767 234 779
rect 200 711 234 729
rect 200 695 234 711
rect 200 643 234 657
rect 200 623 234 643
rect 658 1357 692 1377
rect 658 1343 692 1357
rect 658 1289 692 1305
rect 658 1271 692 1289
rect 658 1221 692 1233
rect 658 1199 692 1221
rect 658 1153 692 1161
rect 658 1127 692 1153
rect 658 1085 692 1089
rect 658 1055 692 1085
rect 658 983 692 1017
rect 658 915 692 945
rect 658 911 692 915
rect 658 847 692 873
rect 658 839 692 847
rect 658 779 692 801
rect 658 767 692 779
rect 658 711 692 729
rect 658 695 692 711
rect 658 643 692 657
rect 658 623 692 643
rect 371 -17 405 17
<< metal1 >>
rect 90 1897 704 1940
rect 90 1863 371 1897
rect 405 1863 704 1897
rect 90 1820 704 1863
rect 194 1377 240 1400
rect 194 1343 200 1377
rect 234 1343 240 1377
rect 194 1305 240 1343
rect 194 1271 200 1305
rect 234 1271 240 1305
rect 194 1233 240 1271
rect 194 1199 200 1233
rect 234 1199 240 1233
rect 194 1161 240 1199
rect 194 1127 200 1161
rect 234 1127 240 1161
rect 194 1089 240 1127
rect 194 1055 200 1089
rect 234 1055 240 1089
rect 194 1017 240 1055
rect 194 983 200 1017
rect 234 983 240 1017
rect 194 945 240 983
rect 194 911 200 945
rect 234 911 240 945
rect 194 873 240 911
rect 194 839 200 873
rect 234 839 240 873
rect 194 801 240 839
rect 194 767 200 801
rect 234 767 240 801
rect 194 729 240 767
rect 194 695 200 729
rect 234 695 240 729
rect 194 657 240 695
rect 194 623 200 657
rect 234 623 240 657
rect 194 600 240 623
rect 652 1377 698 1400
rect 652 1343 658 1377
rect 692 1343 698 1377
rect 652 1305 698 1343
rect 652 1271 658 1305
rect 692 1271 698 1305
rect 652 1233 698 1271
rect 652 1199 658 1233
rect 692 1199 698 1233
rect 652 1161 698 1199
rect 652 1127 658 1161
rect 692 1127 698 1161
rect 652 1089 698 1127
rect 652 1055 658 1089
rect 692 1055 698 1089
rect 652 1017 698 1055
rect 652 983 658 1017
rect 692 983 698 1017
rect 652 945 698 983
rect 652 911 658 945
rect 692 911 698 945
rect 652 873 698 911
rect 652 839 658 873
rect 692 839 698 873
rect 652 801 698 839
rect 652 767 658 801
rect 692 767 698 801
rect 652 729 698 767
rect 652 695 658 729
rect 692 695 698 729
rect 652 657 698 695
rect 652 623 658 657
rect 692 623 698 657
rect 652 600 698 623
rect 90 17 704 60
rect 90 -17 371 17
rect 405 -17 704 17
rect 90 -60 704 -17
<< labels >>
flabel locali s 644 144 704 204 1 FreeSans 1250 0 0 0 GATE
port 1 nsew
flabel locali s 644 1690 704 1750 1 FreeSans 1250 0 0 0 SOURCE
port 2 nsew
flabel locali s 644 370 704 430 1 FreeSans 1250 0 0 0 DRAIN
port 3 nsew
flabel metal1 s 188 1850 248 1910 1 FreeSans 1250 0 0 0 VPWR
port 4 nsew
flabel metal1 s 188 -30 248 30 1 FreeSans 1250 0 0 0 VGND
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 794 1880
<< end >>
