magic
tech sky130A
magscale 1 2
timestamp 1654804491
<< metal3 >>
rect 510520 699926 515374 703728
rect 520526 702378 525364 703622
rect 510508 699688 515374 699926
rect 510508 697518 515372 699688
rect 520502 697586 525388 702378
rect 510520 695072 515372 697518
rect 520526 695031 525364 697586
rect 570344 639766 583336 644534
rect 570508 629776 583360 634544
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0 ~/ee372/caravel_user_project_analog_BGR/mag
timestamp 1632839657
transform 1 0 -46 0 1 -34
box -800 -800 584800 704800
<< labels >>
flabel metal3 572794 639892 580354 644504 1 FreeSans 8000 0 0 0 VCCD1
flabel metal3 510540 698746 515362 701146 1 FreeSans 8000 0 0 0 VSSA1
<< end >>
