magic
tech sky130A
magscale 1 2
timestamp 1654860894
<< metal1 >>
rect 573584 494882 573796 494888
rect 565696 494762 573796 494882
rect 565696 493760 565816 494762
rect 566176 494126 566186 494310
rect 566408 494126 566418 494310
rect 559792 492548 560110 492554
rect 559788 492536 560448 492548
rect 559788 492324 559802 492536
rect 560012 492340 560448 492536
rect 566196 492512 566404 494126
rect 573584 493658 573796 494762
rect 580846 494136 580856 494348
rect 581040 494136 581050 494348
rect 573584 493654 573980 493658
rect 560012 492324 560340 492340
rect 559788 492304 560340 492324
rect 566034 492304 566404 492512
rect 573576 493534 575408 493654
rect 559788 492000 559996 492304
rect 573576 492196 573796 493534
rect 573506 492160 573954 492196
rect 559788 491884 560792 492000
rect 559834 491880 560792 491884
rect 565726 491604 565846 492000
rect 573506 491888 573564 492160
rect 573874 492076 573954 492160
rect 580852 492130 581040 494136
rect 573874 491948 575038 492076
rect 580660 492026 581040 492130
rect 573874 491888 574934 491948
rect 573506 491868 574934 491888
rect 575288 491604 575408 491774
rect 565726 491484 575408 491604
rect 560592 406072 573714 406192
rect 560592 404618 560712 406072
rect 566254 405476 566462 405488
rect 566246 405258 566256 405476
rect 566462 405258 566472 405476
rect 563520 404618 565944 404738
rect 559706 403370 560120 403492
rect 559706 403368 560238 403370
rect 559706 403280 559736 403368
rect 559704 403192 559736 403280
rect 559926 403192 560238 403368
rect 559704 403162 560238 403192
rect 566254 403162 566462 405258
rect 573512 404778 573714 406072
rect 580076 405402 580180 405420
rect 580064 405292 580074 405402
rect 580182 405292 580192 405402
rect 573512 404658 574704 404778
rect 573512 403353 573672 404658
rect 573509 403312 574144 403353
rect 559704 402858 560146 403162
rect 573509 403107 573538 403312
rect 573510 402980 573538 403107
rect 573888 403120 574144 403312
rect 580076 403254 580180 405292
rect 579938 403150 580180 403254
rect 573888 403084 574194 403120
rect 573888 402980 574196 403084
rect 573510 402956 574196 402980
rect 559704 402738 560846 402858
rect 561520 402738 574718 402858
rect 565736 360464 573796 360584
rect 565736 359300 565856 360464
rect 566270 359978 566494 360002
rect 566264 359786 566274 359978
rect 566500 359786 566510 359978
rect 559702 357844 559712 358052
rect 559920 357844 560194 358052
rect 566270 357846 566494 359786
rect 573588 359350 573796 360464
rect 580252 359906 580356 359934
rect 580242 359786 580252 359906
rect 580358 359786 580368 359906
rect 573588 359256 574882 359350
rect 573590 359230 574882 359256
rect 573590 357965 573828 359230
rect 573509 357959 573828 357965
rect 573509 357920 573911 357959
rect 566270 357844 566418 357846
rect 559732 357540 559928 357844
rect 573509 357594 573540 357920
rect 573878 357810 573911 357920
rect 580252 357826 580356 359786
rect 573878 357682 574512 357810
rect 580134 357722 580356 357826
rect 573878 357594 574390 357682
rect 573509 357564 574390 357594
rect 559732 357420 560670 357540
rect 565760 357422 566070 357542
rect 565950 357230 566070 357422
rect 574762 357230 574882 357470
rect 565950 357110 574882 357230
rect 508352 356446 508362 356582
rect 508652 356446 508662 356582
rect 565598 314298 573770 314418
rect 565598 312992 565718 314298
rect 566116 313610 566126 313804
rect 566346 313794 566356 313804
rect 566346 313610 566362 313794
rect 559642 311536 559652 311744
rect 559860 311536 560094 311744
rect 566116 311536 566362 313610
rect 573546 313182 573770 314298
rect 580844 313778 580948 313782
rect 580756 313770 580948 313778
rect 580748 313602 580758 313770
rect 580944 313602 580954 313770
rect 573546 313062 575350 313182
rect 573546 311742 573800 313062
rect 573432 311700 574046 311742
rect 559648 311232 559880 311536
rect 573432 311420 573492 311700
rect 573834 311590 574046 311700
rect 580756 311658 580948 313602
rect 573834 311420 574952 311590
rect 580578 311554 580948 311658
rect 573432 311392 574952 311420
rect 573432 311382 574050 311392
rect 575096 311240 575330 311302
rect 559648 311172 565664 311232
rect 575092 311172 575350 311240
rect 559648 311052 575350 311172
<< via1 >>
rect 566186 494126 566408 494310
rect 559802 492324 560012 492536
rect 580856 494136 581040 494348
rect 573564 491888 573874 492160
rect 566256 405258 566462 405476
rect 559736 403192 559926 403368
rect 580074 405292 580182 405402
rect 573538 402980 573888 403312
rect 566274 359786 566500 359978
rect 559712 357844 559920 358052
rect 580252 359786 580358 359906
rect 573540 357594 573878 357920
rect 508362 356446 508652 356582
rect 566126 313610 566346 313804
rect 559652 311536 559860 311744
rect 580758 313602 580944 313770
rect 573492 311420 573834 311700
<< metal2 >>
rect 580856 494348 581040 494358
rect 566186 494310 566408 494320
rect 580856 494126 581040 494136
rect 566186 494116 566408 494126
rect 559802 492536 560012 492546
rect 559802 492314 560012 492324
rect 573564 492160 573874 492170
rect 573564 491878 573874 491888
rect 566256 405476 566462 405486
rect 580074 405402 580182 405412
rect 580074 405282 580182 405292
rect 566256 405248 566462 405258
rect 559736 403368 559926 403378
rect 559736 403182 559926 403192
rect 573538 403312 573888 403322
rect 573538 402970 573888 402980
rect 541952 389470 542058 389480
rect 541952 389378 542058 389388
rect 541958 380644 542066 380654
rect 542066 380564 542068 380620
rect 541958 380562 542068 380564
rect 541958 380554 542066 380562
rect 566274 359978 566500 359988
rect 566274 359776 566500 359786
rect 580252 359906 580358 359916
rect 580252 359776 580358 359786
rect 559712 358052 559920 358062
rect 559712 357834 559920 357844
rect 573540 357920 573878 357930
rect 573540 357584 573878 357594
rect 508362 356582 508652 356592
rect 508362 356436 508652 356446
rect 566126 313804 566346 313814
rect 566126 313600 566346 313610
rect 580758 313770 580944 313780
rect 580758 313592 580944 313602
rect 559652 311744 559860 311754
rect 559652 311526 559860 311536
rect 573492 311700 573834 311710
rect 573492 311410 573834 311420
<< via2 >>
rect 566186 494126 566408 494310
rect 580856 494136 581040 494348
rect 559802 492324 560012 492536
rect 573564 491888 573874 492160
rect 566256 405258 566462 405476
rect 580074 405292 580182 405402
rect 559736 403192 559926 403368
rect 573538 402980 573888 403312
rect 541952 389388 542058 389470
rect 541958 380564 542066 380644
rect 566274 359786 566500 359978
rect 580252 359786 580358 359906
rect 559712 357844 559920 358052
rect 573540 357594 573878 357920
rect 508362 356446 508652 356582
rect 566126 313610 566346 313804
rect 580758 313602 580944 313770
rect 559652 311536 559860 311744
rect 573492 311420 573834 311700
<< metal3 >>
rect 413300 698232 418436 703282
rect 465296 698476 470432 703526
rect 510560 701276 515394 703604
rect 510552 701180 515394 701276
rect 510552 700092 515386 701180
rect 510552 699264 515392 700092
rect 510538 697668 515392 699264
rect 510538 697378 515372 697668
rect 510538 696840 510704 697378
rect 510560 689882 510704 696840
rect 515202 689882 515372 697378
rect 510560 689666 515372 689882
rect 520554 697354 525388 703122
rect 566500 698354 571636 703404
rect 520554 689858 520704 697354
rect 525202 689858 525388 697354
rect 520554 689727 525388 689858
rect 577256 677954 582392 683004
rect 567105 644596 581232 644606
rect 567105 644324 582918 644596
rect 567105 640080 567306 644324
rect 573722 640080 582918 644324
rect 567105 639760 582918 640080
rect 567308 634256 583176 634588
rect 567296 630012 567306 634256
rect 573722 630012 583176 634256
rect 567308 629752 583176 630012
rect 580846 494348 581050 494353
rect 566148 494310 566454 494332
rect 566148 494248 566186 494310
rect 501828 494126 566186 494248
rect 566408 494248 566454 494310
rect 580846 494248 580856 494348
rect 566408 494136 580856 494248
rect 581040 494248 581050 494348
rect 581040 494136 583862 494248
rect 566408 494126 583862 494136
rect 501828 494124 583862 494126
rect 501828 415012 501952 494124
rect 566148 494090 566454 494124
rect 559792 492536 560022 492541
rect 559792 492324 559802 492536
rect 560012 492324 560022 492536
rect 559792 492319 560022 492324
rect 573554 492160 573884 492165
rect 573554 491888 573564 492160
rect 573874 491888 573884 492160
rect 573554 491883 573884 491888
rect 501026 414806 501952 415012
rect 566246 405476 566472 405481
rect 566246 405400 566256 405476
rect 542962 405288 566256 405400
rect 542962 389490 543074 405288
rect 566246 405258 566256 405288
rect 566462 405400 566472 405476
rect 580064 405402 580192 405407
rect 580064 405400 580074 405402
rect 566462 405292 580074 405400
rect 580182 405400 580192 405402
rect 580182 405292 583872 405400
rect 566462 405288 583872 405292
rect 566462 405258 566472 405288
rect 580064 405287 580192 405288
rect 566246 405253 566472 405258
rect 559726 403368 559936 403373
rect 559726 403192 559736 403368
rect 559926 403192 559936 403368
rect 559726 403187 559936 403192
rect 573528 403312 573898 403317
rect 573528 402980 573538 403312
rect 573888 402980 573898 403312
rect 573528 402975 573898 402980
rect 541910 389470 543074 389490
rect 541910 389388 541952 389470
rect 542058 389388 543074 389470
rect 541910 389378 543074 389388
rect 541937 380644 545137 380703
rect 541937 380564 541958 380644
rect 542066 380615 545137 380644
rect 542066 380564 545141 380615
rect 541937 380499 545141 380564
rect 541959 380497 545141 380499
rect 545023 359903 545141 380497
rect 566264 359978 566510 359983
rect 566264 359903 566274 359978
rect 545023 359786 566274 359903
rect 566500 359903 566510 359978
rect 580242 359906 580368 359911
rect 580242 359903 580252 359906
rect 566500 359786 580252 359903
rect 580358 359903 580368 359906
rect 580358 359786 580941 359903
rect 545023 359785 580941 359786
rect 566264 359781 566510 359785
rect 580242 359781 580368 359785
rect 580823 358984 580941 359785
rect 580823 358866 583840 358984
rect 580823 358859 580941 358866
rect 559702 358052 559930 358057
rect 559702 357844 559712 358052
rect 559920 357844 559930 358052
rect 559702 357839 559930 357844
rect 573530 357920 573888 357925
rect 573530 357594 573540 357920
rect 573878 357594 573888 357920
rect 573530 357589 573888 357594
rect 508335 356582 509603 356589
rect 508335 356446 508362 356582
rect 508652 356446 509603 356582
rect 508335 356375 509603 356446
rect 509393 313770 509603 356375
rect 566116 313804 566356 313809
rect 566116 313770 566126 313804
rect 509393 313610 566126 313770
rect 566346 313770 566356 313804
rect 580748 313770 580954 313775
rect 566346 313610 580758 313770
rect 509393 313602 580758 313610
rect 580944 313727 583738 313770
rect 580944 313602 583873 313727
rect 509393 313593 583873 313602
rect 559642 311744 559870 311749
rect 559642 311536 559652 311744
rect 559860 311536 559870 311744
rect 559642 311531 559870 311536
rect 573482 311700 573844 311705
rect 573482 311420 573492 311700
rect 573834 311420 573844 311700
rect 573482 311415 573844 311420
<< via3 >>
rect 510704 689882 515202 697378
rect 520704 689858 525202 697354
rect 567306 640080 573722 644324
rect 567306 630012 573722 634256
rect 559802 492324 560012 492536
rect 573564 491888 573874 492160
rect 559736 403192 559926 403368
rect 573538 402980 573888 403312
rect 559712 357844 559920 358052
rect 573540 357594 573878 357920
rect 559652 311536 559860 311744
rect 573492 311420 573834 311700
<< metal4 >>
rect 502376 697378 560022 697790
rect 502376 689882 510704 697378
rect 515202 697354 560022 697378
rect 515202 689882 520704 697354
rect 502376 689858 520704 689882
rect 525202 689858 560022 697354
rect 502376 689742 560022 689858
rect 551974 492536 560022 689742
rect 567305 644324 573723 644325
rect 567305 640080 567306 644324
rect 573722 640080 573723 644324
rect 567305 640079 573723 640080
rect 567305 634256 573723 634257
rect 567305 630012 567306 634256
rect 573722 630012 573723 634256
rect 567305 630011 573723 630012
rect 551974 492324 559802 492536
rect 560012 492324 560022 492536
rect 551974 414054 560022 492324
rect 573563 492160 573875 492161
rect 573563 491888 573564 492160
rect 573874 491888 573875 492160
rect 573563 491887 573875 491888
rect 529718 412422 560022 414054
rect 551974 403368 560022 412422
rect 551974 403192 559736 403368
rect 559926 403192 560022 403368
rect 551974 359050 560022 403192
rect 573537 403312 573889 403313
rect 573537 402980 573538 403312
rect 573888 402980 573889 403312
rect 573537 402979 573889 402980
rect 528872 358052 560022 359050
rect 528872 357844 559712 358052
rect 559920 357844 560022 358052
rect 528872 357418 560022 357844
rect 573539 357920 573879 357921
rect 573539 357594 573540 357920
rect 573878 357594 573879 357920
rect 573539 357593 573879 357594
rect 551974 311744 560022 357418
rect 551974 311536 559652 311744
rect 559860 311536 560022 311744
rect 551974 154934 560022 311536
rect 573491 311700 573835 311701
rect 573491 311420 573492 311700
rect 573834 311420 573835 311700
rect 573491 311419 573835 311420
<< via4 >>
rect 567306 640080 573722 644324
rect 567306 630012 573722 634256
rect 573564 491888 573874 492160
rect 573538 402980 573888 403312
rect 573540 357594 573878 357920
rect 573492 311420 573834 311700
<< metal5 >>
rect 567158 644324 573920 649062
rect 567158 640080 567306 644324
rect 573722 640080 573920 644324
rect 567158 634256 573920 640080
rect 567158 630012 567306 634256
rect 573722 630012 573920 634256
rect 567158 627314 573920 630012
rect 567156 621952 573942 627314
rect 567158 492160 573920 621952
rect 567158 491888 573564 492160
rect 573874 491888 573920 492160
rect 488780 422974 490412 423442
rect 567158 422974 573920 491888
rect 488780 421342 573920 422974
rect 488780 405016 490412 421342
rect 536984 420968 573920 421342
rect 537164 401694 538796 420968
rect 567158 403312 573920 420968
rect 567158 402980 573538 403312
rect 573888 402980 573920 403312
rect 488780 348924 490412 365430
rect 537164 348924 538796 366466
rect 567158 357920 573920 402980
rect 567158 357594 573540 357920
rect 573878 357594 573920 357920
rect 567158 348924 573920 357594
rect 488668 347292 573920 348924
rect 567158 311700 573920 347292
rect 567158 311420 573492 311700
rect 573834 311420 573920 311700
rect 567158 147385 573920 311420
use bgr_top_flat  bgr_top_flat_0 ~/ee372/caravel_user_project_analog_BGR/mag
timestamp 1654805184
transform 0 -1 542060 -1 0 414954
box 0 0 58516 56576
use nmos_flat  nmos_flat_0
timestamp 1654813604
transform -1 0 563258 0 1 492940
box -3268 -1060 3164 940
use nmos_flat  nmos_flat_1
timestamp 1654813604
transform -1 0 563194 0 1 403798
box -3268 -1060 3164 940
use nmos_flat  nmos_flat_2
timestamp 1654813604
transform -1 0 563150 0 1 358480
box -3268 -1060 3164 940
use nmos_flat  nmos_flat_3
timestamp 1654813604
transform -1 0 563012 0 1 312172
box -3268 -1060 3164 940
use pmos_flat  pmos_flat_0
timestamp 1654850744
transform -1 0 577092 0 1 403838
box -2950 -1060 3026 940
use pmos_flat  pmos_flat_1
timestamp 1654850744
transform -1 0 577288 0 1 358410
box -2950 -1060 3026 940
use pmos_flat  pmos_flat_2
timestamp 1654850744
transform -1 0 577736 0 1 312242
box -2950 -1060 3026 940
use pmos_flat  pmos_flat_3
timestamp 1654850744
transform -1 0 577814 0 1 492714
box -2950 -1060 3026 940
use user_analog_project_wrapper_empty  user_analog_project_wrapper_empty_0
timestamp 1632839657
transform 1 0 -24 0 1 -12
box -800 -800 584800 704800
<< labels >>
flabel metal3 510596 697782 515352 701406 1 FreeSans 8000 0 0 0 VSSA1
flabel metal3 574704 639800 581232 644606 1 FreeSans 8000 0 0 0 VCCD1
<< end >>
