magic
tech sky130A
timestamp 1655503347
<< metal4 >>
rect -408 379 408 408
rect -408 -379 -379 379
rect 379 -379 408 379
rect -408 -408 408 -379
<< via4 >>
rect -379 -379 379 379
<< metal5 >>
rect -408 379 408 408
rect -408 -379 -379 379
rect 379 -379 408 379
rect -408 -408 408 -379
<< end >>
