* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt bgr_all_flat nmos_flat_3/VPWR pmos_flat_2/VGND bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rout
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/Rin bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/Rin
+ bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/Rin bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE
+ bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN nmos_flat_0/VPWR
+ nmos_flat_1/VPWR nmos_flat_2/VPWR VSSA1 pmos_flat_0/VGND nmos_flat_1/GATE pmos_flat_1/VGND
+ pmos_flat_1/DRAIN pmos_flat_3/VGND pmos_flat_3/DRAIN VCCD1 m3_413300_698232# pmos_flat_1/VPWR
+ m3_566500_698354# pmos_flat_2/VPWR pmos_flat_3/VPWR m3_465296_698476# pmos_flat_0/VPWR
+ m3_577256_677954#
X0 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=3.2244e+14p pd=1.90726e+09u as=1.45e+13p ps=1.058e+08u w=5e+06u l=1e+06u
X1 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+13p ps=1.058e+08u w=5e+06u l=1e+06u
X2 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X3 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=2.60014e+14p pd=1.87904e+09u as=7.39355e+13p ps=5.3426e+08u w=6.45e+06u l=2e+06u
X4 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+13p ps=1.058e+08u w=5e+06u l=1e+06u
X5 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X7 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=9.8589e+13p pd=6.4222e+08u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 VSSA1 VSSA1 a_560541_357980# VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X10 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X11 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 a_515903_369632# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X13 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X14 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=1.45e+13p pd=1.058e+08u as=0p ps=0u w=5e+06u l=1e+06u
X15 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X16 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X17 a_565849_403298# nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=1e+06u
X18 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X20 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=7.39355e+13p pd=5.3426e+08u as=0p ps=0u w=6.45e+06u l=2e+06u
X21 a_519663_379334# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X22 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X23 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X24 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X25 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X26 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X27 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X28 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X29 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X30 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X31 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X32 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X33 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X34 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X35 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X36 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X37 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X38 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X39 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X40 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X41 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X42 a_519663_388644# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X43 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X44 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.30935e+13p ps=9.436e+07u w=6.45e+06u l=2e+06u
X45 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X46 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X47 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X48 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X49 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X50 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X51 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X52 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X53 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X54 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.595e+13p ps=1.1638e+08u w=5e+06u l=1e+06u
X55 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X56 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X57 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X58 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X59 a_493343_391682# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X60 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X61 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X62 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X63 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X64 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X65 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X66 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X67 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X68 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X69 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X70 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X71 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X72 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X73 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X74 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X75 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X76 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X77 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X78 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X79 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X80 a_530943_368750# pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X81 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X82 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X83 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X84 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X85 a_515903_390114# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X86 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X87 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X88 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X89 a_519663_385312# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X90 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X91 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X92 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=1.16e+13p pd=8.58e+07u as=0p ps=0u w=4e+06u l=2e+06u
X93 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X94 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X95 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X96 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X97 VSSA1 nmos_flat_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X98 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X99 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X100 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X101 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X102 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X103 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X104 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X105 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.276e+13p ps=9.438e+07u w=4e+06u l=2e+06u
X106 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X107 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X108 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X109 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X110 a_530943_363262# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X111 a_504623_390016# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X112 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X113 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X114 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X115 a_504623_398836# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X116 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X117 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X118 a_534703_367966# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X119 VCCD1 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=7.482e+12p ps=5.392e+07u w=6.45e+06u l=2e+06u
X120 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X121 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X122 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X123 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X124 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X125 a_519663_364144# pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X126 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X127 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X128 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X129 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X130 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X131 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X133 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X134 a_504623_392773# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X135 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X136 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X137 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X138 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X139 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X140 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X141 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X142 a_512143_393250# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X143 a_504623_396092# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X144 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X145 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X146 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X147 a_534703_365222# VSSA1 VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X148 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X149 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X150 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X151 a_519663_382568# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X152 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X153 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X154 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X155 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X156 VCCD1 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X157 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X158 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X159 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X160 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X161 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X162 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X163 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X164 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X165 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X166 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X167 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X169 a_515903_375120# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X170 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X171 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X172 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X173 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X174 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X175 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X176 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X177 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X178 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X179 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X180 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X181 a_534703_362478# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X182 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X183 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X184 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X185 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=5.8e+12p pd=4.29e+07u as=0p ps=0u w=4e+06u l=2e+06u
X186 VCCD1 VCCD1 pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X187 a_527183_368652# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X188 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X189 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X190 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X191 a_519663_385312# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rout VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X192 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X193 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X194 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X195 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X196 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X197 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X198 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X199 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X200 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X201 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X202 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X203 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X204 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X206 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X207 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X208 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X209 a_527183_363164# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X210 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X211 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X212 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X213 VCCD1 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=7.482e+12p ps=5.392e+07u w=6.45e+06u l=2e+06u
X214 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X215 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X216 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X217 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X218 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X219 a_527183_365908# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X220 a_519663_372376# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X221 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X222 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=2e+06u
X223 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X224 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X225 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X226 pmos_flat_3/DRAIN VCCD1 VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X227 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X228 a_515903_369632# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X229 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X230 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X231 a_519663_364144# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X232 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X233 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X234 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X235 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X236 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X237 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X238 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X239 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X240 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X241 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X242 a_512143_395994# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X243 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X244 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X245 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X246 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X247 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X248 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X249 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X250 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X251 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X252 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X253 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X254 a_508383_389931# VSSA1 VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X255 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X256 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X257 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X258 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X259 VCCD1 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X260 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X261 VSSA1 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__pnp_05v5 area=0p
X262 a_519663_382568# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X263 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X264 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X265 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X266 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X267 a_508383_393250# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X268 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X269 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X270 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X271 a_512143_390506# pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X272 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X273 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X274 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X275 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X276 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X277 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X278 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X279 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X280 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X281 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X282 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X283 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X284 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X285 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X286 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X287 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X288 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X289 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X290 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X291 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X292 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X293 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X294 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X295 a_530943_366006# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X296 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X297 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X298 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X299 a_515903_390114# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X300 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X301 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X302 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X303 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X304 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X305 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X306 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X307 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X308 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X309 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X310 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X311 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X312 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X313 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X314 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X315 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X316 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X317 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X318 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X319 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X320 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X321 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X322 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X323 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X324 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X325 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X326 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X327 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X328 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X329 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X330 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X331 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X332 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X333 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X334 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X335 VCCD1 VCCD1 pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X336 a_504623_390016# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X337 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X338 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X339 VCCD1 VCCD1 pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X340 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X341 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X342 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X343 a_534703_367966# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X344 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X345 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X346 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X347 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X348 a_519663_372376# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X349 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X350 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X351 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X352 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X353 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X354 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X355 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X356 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X357 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X358 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X359 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X360 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X361 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X362 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X363 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X364 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X365 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X366 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X367 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X368 a_493343_391682# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X369 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X370 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X371 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X372 a_515903_364144# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X373 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X374 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X375 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X376 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X377 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X378 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X379 VCCD1 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X380 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X381 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X382 a_515903_366888# pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X383 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X384 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X385 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X386 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X387 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X388 a_534703_365222# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X389 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X390 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X391 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X392 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X393 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X394 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X395 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X396 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X397 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X398 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X399 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X400 a_512143_385312# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X401 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X402 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X403 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X404 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X405 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X406 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X407 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X408 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X409 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X410 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X411 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X412 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X413 a_519663_375120# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X414 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X415 VCCD1 VCCD1 pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X416 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X417 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X418 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X419 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X420 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X421 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X422 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X423 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X424 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X425 a_534703_362478# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X426 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X427 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X428 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X429 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X430 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X431 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X432 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X433 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X434 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X435 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X436 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X437 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X438 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X439 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X440 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X441 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X442 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X443 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X444 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X445 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X446 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X447 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X448 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X449 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X450 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X451 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X452 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X453 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X454 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X455 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X456 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X457 pmos_flat_3/DRAIN VCCD1 VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X458 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X459 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X460 pmos_flat_3/DRAIN VCCD1 VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X461 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X462 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X463 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X464 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X465 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X466 a_512143_393250# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X467 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X468 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X469 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X470 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X471 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X472 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X473 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X474 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X475 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X476 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X477 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X478 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X479 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X480 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X481 VSSA1 VSSA1 a_560403_311672# VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X482 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X483 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X484 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X485 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X486 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X487 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X488 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X489 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X490 a_515903_372376# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X491 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X492 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X493 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X494 VSSA1 VSSA1 a_560649_492440# VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u l=1e+06u
X495 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X496 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X497 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X498 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X499 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X500 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X501 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X502 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X503 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X504 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X505 a_530943_368750# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X506 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X507 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X508 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X509 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X510 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X511 VCCD1 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X512 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X513 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X514 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X515 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X516 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X517 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X518 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X519 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X520 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X521 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X522 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X523 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X524 a_527183_368652# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X525 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X526 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X527 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X528 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X529 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X530 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X531 a_530943_363262# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X532 pmos_flat_3/DRAIN VCCD1 VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X533 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X534 pmos_flat_3/DRAIN VCCD1 VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X535 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X536 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X537 a_519663_375120# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X538 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X539 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X540 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X541 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X542 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X543 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X544 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X545 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X546 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X547 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X548 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X549 a_527183_363164# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X550 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X551 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X552 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X553 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X554 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X555 a_527183_365908# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X556 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X557 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X558 VSSA1 nmos_flat_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X559 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X560 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X561 VSSA1 nmos_flat_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X562 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X563 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X564 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X565 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X566 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X567 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X568 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X569 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X570 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X571 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X572 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X573 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X574 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X575 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X576 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X577 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X578 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X579 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X580 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X581 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X582 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X583 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X584 VSSA1 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X585 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X586 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X587 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X588 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X589 a_508383_389931# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X590 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X591 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X592 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X593 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X594 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X595 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X596 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X597 a_508383_393250# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X598 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X599 VSSA1 nmos_flat_1/GATE bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X600 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X601 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X602 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X603 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X604 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X605 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X606 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X607 pmos_flat_1/DRAIN VCCD1 VCCD1 pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X608 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X609 a_504623_398836# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X610 a_515903_364144# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X611 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X612 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X613 a_515903_366888# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X614 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X615 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X616 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X617 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X618 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X619 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X620 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X621 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X622 VCCD1 VCCD1 nmos_flat_1/GATE pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X623 a_530943_366006# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X624 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X625 a_519663_379334# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X626 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X627 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X628 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X629 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X630 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X631 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X632 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X633 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X634 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X635 a_504623_392773# VSSA1 VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X636 VCCD1 VCCD1 pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X637 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X638 VCCD1 VCCD1 pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X639 bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X640 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X641 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X642 pmos_flat_2/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X643 pmos_flat_3/DRAIN VCCD1 VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X644 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X645 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X646 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X647 a_504623_396092# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X648 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X649 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X650 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X651 pmos_flat_3/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X652 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X653 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X654 a_519663_388644# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X655 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X656 pmos_flat_3/DRAIN VCCD1 VCCD1 pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X657 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X658 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X659 VSSA1 VSSA1 pmos_flat_1/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X660 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X661 VSSA1 VSSA1 pmos_flat_3/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X662 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X663 VSSA1 VSSA1 bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_fd_pr__pnp_05v5 area=0p
X664 VCCD1 VCCD1 pmos_flat_3/DRAIN pmos_flat_3/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X665 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X666 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X667 pmos_flat_1/DRAIN VSSA1 VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X668 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X669 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X670 nmos_flat_1/GATE nmos_flat_1/GATE VSSA1 VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X671 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X672 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X673 a_515903_375120# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X674 a_512143_395994# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X675 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X676 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X677 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X678 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X679 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X680 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X681 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X682 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_2/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X683 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X684 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X685 bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X686 VCCD1 VCCD1 pmos_flat_1/DRAIN pmos_flat_1/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X687 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X688 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X689 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X690 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_3/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X691 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X692 VSSA1 pmos_flat_3/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X693 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X694 pmos_flat_3/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X695 a_512143_390506# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X696 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X697 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X698 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X699 pmos_flat_2/DRAIN VCCD1 VCCD1 pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X700 VCCD1 VCCD1 pmos_flat_2/DRAIN pmos_flat_2/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X701 pmos_flat_1/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X702 nmos_flat_1/GATE VCCD1 VCCD1 pmos_flat_0/VPWR sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X703 VSSA1 VSSA1 pmos_flat_2/DRAIN VSSA1 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X704 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X705 VCCD1 bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout pmos_flat_1/DRAIN VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X706 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X707 a_512143_385312# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rout VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X708 a_515903_372376# bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/Rin VSSA1 sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X709 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X710 pmos_flat_2/DRAIN bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout VCCD1 VCCD1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[4] io_analog[5] io_analog[6] io_analog[7]
+ io_analog[8] io_analog[9] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
Xbgr_all_flat_0 bgr_all_flat_0/nmos_flat_3/VPWR bgr_all_flat_0/pmos_flat_2/VGND bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_1/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_2/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_4/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_6/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_7/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_5/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_8/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_0/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_12/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_10/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_19/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_13/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_18/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_17/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_11/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_20/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_24/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_23/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_9/Rout
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_0/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_16/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_28/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_27/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_29/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_2_1/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_pfet_01v8_lvt_6_1/GATE bgr_all_flat_0/bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_0/DRAIN
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_21/Rout bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_30/Rin
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_res_xhigh_po_2p85_1_26/Rin bgr_all_flat_0/bgr_top_flat_0/sky130_asc_nfet_01v8_lvt_1_1/GATE
+ bgr_all_flat_0/bgr_top_flat_0/sky130_asc_cap_mim_m3_1_4/Cout gpio_analog[1] bgr_all_flat_0/nmos_flat_0/VPWR
+ bgr_all_flat_0/nmos_flat_1/VPWR bgr_all_flat_0/nmos_flat_2/VPWR vssa1 bgr_all_flat_0/pmos_flat_0/VGND
+ gpio_analog[3] bgr_all_flat_0/pmos_flat_1/VGND gpio_analog[2] bgr_all_flat_0/pmos_flat_3/VGND
+ gpio_analog[5] vccd1 io_analog[3] bgr_all_flat_0/pmos_flat_1/VPWR io_analog[1] bgr_all_flat_0/pmos_flat_2/VPWR
+ bgr_all_flat_0/pmos_flat_3/VPWR io_analog[2] bgr_all_flat_0/pmos_flat_0/VPWR io_analog[0]
+ bgr_all_flat
.ends

