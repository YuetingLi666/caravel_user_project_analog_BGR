magic
tech sky130A
magscale 1 2
timestamp 1655764969
<< locali >>
rect 423954 689608 424312 689668
rect 406576 689458 406890 689498
rect 406636 687976 406676 689458
rect 418324 688288 418906 688348
rect 424252 688202 424312 689608
rect 458334 689644 458742 689660
rect 458266 689620 458742 689644
rect 458266 689584 458390 689620
rect 411986 688078 413262 688138
rect 423904 688122 424234 688182
rect 458330 688138 458390 689584
rect 476236 689574 476642 689634
rect 463788 688240 465158 688300
rect 470670 688254 471182 688314
rect 476582 688184 476642 689574
rect 458330 688078 458758 688138
rect 476292 688088 476550 688148
rect 406636 687916 407198 687976
rect 560520 582856 560827 582916
rect 560520 581430 560580 582856
rect 574316 582752 574638 582792
rect 565923 581536 566340 581596
rect 560362 581428 560908 581430
rect 560406 581370 560908 581428
rect 574316 581270 574356 582752
rect 579714 581372 580148 581432
rect 574344 581210 574746 581270
rect 574532 509262 574850 509302
rect 560374 509174 560758 509234
rect 560374 507764 560434 509174
rect 565840 507854 566212 507914
rect 574532 507800 574572 509262
rect 579986 507882 580388 507942
rect 560450 507686 560782 507746
rect 574586 507720 575030 507780
rect 560392 449212 560622 449272
rect 560392 448050 560452 449212
rect 560288 447990 560452 448050
rect 574700 449018 574960 449058
rect 560392 447784 560452 447990
rect 565715 447898 566266 447952
rect 565715 447892 566364 447898
rect 560392 447724 560624 447784
rect 574700 447534 574740 449018
rect 580050 447638 580686 447698
rect 574428 447478 574889 447534
rect 574303 447476 574889 447478
rect 574388 404536 574676 404576
rect 560374 404224 560704 404284
rect 560374 402798 560434 404224
rect 566392 402964 566452 403310
rect 574388 403054 574428 404536
rect 579754 403156 580108 403216
rect 574327 402994 574740 403054
rect 574388 402990 574428 402994
rect 565749 402904 566452 402964
rect 560270 402738 560726 402798
rect 574432 359110 574696 359150
rect 560398 358756 560620 358816
rect 560186 357426 560208 357518
rect 560148 357328 560208 357426
rect 560398 357328 560458 358756
rect 565676 357438 566298 357496
rect 574432 357628 574472 359110
rect 579802 357730 580280 357790
rect 574332 357570 575022 357628
rect 574196 357568 575022 357570
rect 566444 357438 566454 357496
rect 565676 357436 566454 357438
rect 560148 357268 560570 357328
rect 574840 313042 575074 313082
rect 560306 312820 560654 312880
rect 560306 311680 560366 312820
rect 560246 311620 560366 311680
rect 560306 311394 560366 311620
rect 565606 311508 566156 311560
rect 566358 311508 566380 311560
rect 565606 311500 566380 311508
rect 574840 311560 574880 313042
rect 580246 311662 580536 311722
rect 574718 311500 575232 311560
rect 560306 311334 560826 311394
<< viali >>
rect 406474 689426 406576 689524
rect 418238 688270 418324 688362
rect 458146 689552 458266 689692
rect 413262 688056 413364 688162
rect 424234 688104 424342 688202
rect 465158 688228 465252 688344
rect 470582 688236 470670 688336
rect 476550 688050 476688 688184
rect 566340 581520 566460 581634
rect 560334 581362 560406 581428
rect 580148 581372 580208 581432
rect 574284 581210 574344 581270
rect 566212 507840 566310 507940
rect 580388 507856 580498 507968
rect 560362 507684 560450 507764
rect 574502 507710 574586 507800
rect 560158 447958 560288 448084
rect 566266 447898 566376 448006
rect 574266 447478 574428 447656
rect 580686 447552 580874 447740
rect 560134 402714 560270 402872
rect 566312 403310 566460 403428
rect 574086 402972 574327 403213
rect 580108 403136 580258 403288
rect 560070 357426 560186 357542
rect 566298 357438 566444 357578
rect 574116 357570 574332 357806
rect 580280 357714 580448 357900
rect 560056 311568 560246 311726
rect 566156 311508 566358 311694
rect 574558 311410 574718 311574
rect 580536 311610 580786 311816
<< metal1 >>
rect 423942 691338 424062 691366
rect 423862 691084 423872 691338
rect 424132 691084 424142 691338
rect 476068 691094 476078 691356
rect 476352 691094 476362 691356
rect 423942 689738 424062 691084
rect 458148 689750 458804 689870
rect 406456 689588 407046 689708
rect 458148 689704 458268 689750
rect 476162 689704 476282 691094
rect 458140 689692 458272 689704
rect 406456 689530 406576 689588
rect 458136 689552 458146 689692
rect 458266 689552 458276 689692
rect 458140 689540 458272 689552
rect 406456 689524 406588 689530
rect 406456 689426 406474 689524
rect 406576 689426 406588 689524
rect 406456 689422 406588 689426
rect 406462 689420 406588 689422
rect 418232 688362 418330 688374
rect 418228 688270 418238 688362
rect 418324 688270 418334 688362
rect 465152 688344 465258 688356
rect 418232 688258 418330 688270
rect 465148 688228 465158 688344
rect 465252 688228 465262 688344
rect 470576 688336 470676 688348
rect 470572 688236 470582 688336
rect 470670 688236 470680 688336
rect 465152 688216 465258 688228
rect 470576 688224 470676 688236
rect 424222 688202 424354 688208
rect 413256 688162 413370 688174
rect 413252 688056 413262 688162
rect 413364 688056 413374 688162
rect 424222 688104 424234 688202
rect 424342 688104 424354 688202
rect 424222 688098 424354 688104
rect 476538 688188 476700 688190
rect 476538 688184 476702 688188
rect 413256 688044 413370 688056
rect 424232 687978 424352 688098
rect 476538 688050 476550 688184
rect 476688 688050 476702 688184
rect 476538 688044 476702 688050
rect 423928 687858 424352 687978
rect 463780 687870 464130 687990
rect 476582 687944 476702 688044
rect 412038 686552 412158 687828
rect 412012 686420 412022 686552
rect 412170 686420 412180 686552
rect 464010 686542 464130 687870
rect 476210 687824 476702 687944
rect 463980 686390 463990 686542
rect 464154 686390 464164 686542
rect 464010 686384 464130 686390
rect 437506 668808 437516 668962
rect 437660 668808 437670 668962
rect 446346 668822 446356 668974
rect 446500 668822 446510 668974
rect 565961 583972 574678 584092
rect 565961 582986 566081 583972
rect 566334 583690 566510 583696
rect 566330 583578 566340 583690
rect 566492 583578 566510 583690
rect 566334 581640 566510 583578
rect 574558 583286 574678 583972
rect 580122 583568 580132 583676
rect 580222 583568 580232 583676
rect 566328 581634 566510 581640
rect 559778 581318 559788 581528
rect 560010 581442 560020 581528
rect 566328 581520 566340 581634
rect 566460 581520 566510 581634
rect 566328 581514 566510 581520
rect 573650 583166 574678 583286
rect 560010 581428 560420 581442
rect 573650 581438 573770 583166
rect 574558 582918 574678 583166
rect 580132 581438 580216 583568
rect 560010 581362 560334 581428
rect 560406 581362 560420 581428
rect 560010 581360 560420 581362
rect 560010 581318 560020 581360
rect 560322 581356 560418 581360
rect 559852 581226 559972 581318
rect 559852 581106 560887 581226
rect 565822 581106 572612 581226
rect 573618 581122 573628 581438
rect 573910 581278 573920 581438
rect 580132 581432 580220 581438
rect 580132 581372 580148 581432
rect 580208 581372 580220 581432
rect 580132 581366 580220 581372
rect 573910 581276 574352 581278
rect 573910 581270 574356 581276
rect 573910 581210 574284 581270
rect 574344 581210 574356 581270
rect 573910 581204 574356 581210
rect 573910 581186 574352 581204
rect 573910 581122 573920 581186
rect 572492 580962 572612 581106
rect 574882 580962 575002 581072
rect 572492 580842 575002 580962
rect 574066 509470 574886 509590
rect 574066 509424 574186 509470
rect 565728 509304 574186 509424
rect 566200 507830 566210 507952
rect 566316 507830 566326 507952
rect 573642 507912 573762 509304
rect 580382 507968 580504 507980
rect 566206 507828 566316 507830
rect 559794 507792 559914 507796
rect 559784 507678 559794 507792
rect 559918 507788 559928 507792
rect 559918 507770 560458 507788
rect 559918 507764 560462 507770
rect 559918 507684 560362 507764
rect 560450 507684 560462 507764
rect 559918 507678 560462 507684
rect 559794 507544 559914 507678
rect 573606 507620 573616 507912
rect 573914 507822 573924 507912
rect 580378 507856 580388 507968
rect 580498 507856 580508 507968
rect 580382 507844 580504 507856
rect 573914 507800 574594 507822
rect 573914 507710 574502 507800
rect 574586 507710 574594 507800
rect 573914 507698 574594 507710
rect 573914 507620 573924 507698
rect 559794 507424 560894 507544
rect 565574 507424 573414 507544
rect 573294 507384 573414 507424
rect 574796 507384 574916 507608
rect 573294 507264 574916 507384
rect 573574 450479 573786 450485
rect 565686 450359 573786 450479
rect 565686 449382 565806 450359
rect 566166 449905 566408 449907
rect 566166 449725 566197 449905
rect 566377 449725 566408 449905
rect 566166 449723 566408 449725
rect 566186 449610 566394 449723
rect 559782 448145 560100 448151
rect 559778 448117 560220 448145
rect 559778 447937 559807 448117
rect 559987 448090 560220 448117
rect 559987 448084 560300 448090
rect 559987 447958 560158 448084
rect 560288 447958 560300 448084
rect 566261 448012 566376 449610
rect 573574 449255 573786 450359
rect 580836 449929 581040 449945
rect 580836 449749 580848 449929
rect 581028 449749 581040 449929
rect 580836 449733 581040 449749
rect 574310 449266 574854 449372
rect 573574 449251 573970 449255
rect 574298 449251 574854 449266
rect 573566 449146 574854 449251
rect 573566 449131 574432 449146
rect 559987 447952 560300 447958
rect 566254 448006 566388 448012
rect 559987 447937 560220 447952
rect 559778 447901 560220 447937
rect 559778 447597 559986 447901
rect 566254 447898 566266 448006
rect 566376 447898 566388 448006
rect 566254 447892 566388 447898
rect 573566 447793 573786 449131
rect 573496 447743 573944 447793
rect 580842 447746 581030 449733
rect 559778 447481 560794 447597
rect 559824 447477 560794 447481
rect 565820 447201 565940 447574
rect 573496 447499 573555 447743
rect 573863 447673 573944 447743
rect 580674 447740 581030 447746
rect 573863 447668 574432 447673
rect 573863 447656 574434 447668
rect 573863 447499 574266 447656
rect 573496 447478 574266 447499
rect 574428 447478 574434 447656
rect 580674 447552 580686 447740
rect 580874 447552 581030 447740
rect 580674 447546 580886 447552
rect 573496 447466 574434 447478
rect 573496 447465 574432 447466
rect 574750 447201 574870 447368
rect 565820 447081 574870 447201
rect 560606 406081 573728 406201
rect 560606 404448 560726 406081
rect 566268 405485 566476 405497
rect 566260 405466 566486 405485
rect 566260 405286 566283 405466
rect 566463 405286 566486 405466
rect 566260 405267 566486 405286
rect 566268 405112 566476 405267
rect 559720 403347 559996 403501
rect 566302 403434 566476 405112
rect 559720 403289 559755 403347
rect 559718 403231 559755 403289
rect 559935 403231 559996 403347
rect 566300 403428 566476 403434
rect 566300 403310 566312 403428
rect 566460 403386 566476 403428
rect 573526 404787 573728 406081
rect 580090 405411 580194 405429
rect 580078 405382 580206 405411
rect 580078 405330 580116 405382
rect 580168 405330 580206 405382
rect 580078 405301 580206 405330
rect 574002 404787 574718 404892
rect 573526 404772 574718 404787
rect 573526 404667 574122 404772
rect 566460 403310 566472 403386
rect 573526 403362 573686 404667
rect 566300 403304 566472 403310
rect 573523 403360 574122 403362
rect 573523 403309 574346 403360
rect 559718 403122 559996 403231
rect 559718 402974 560276 403122
rect 573523 403116 573573 403309
rect 560128 402872 560276 402974
rect 573524 403001 573573 403116
rect 573881 403213 574346 403309
rect 573881 403001 574086 403213
rect 573524 402972 574086 403001
rect 574327 402984 574346 403213
rect 580090 403326 580194 405301
rect 580090 403288 580272 403326
rect 580090 403136 580108 403288
rect 580258 403136 580272 403288
rect 580090 403116 580272 403136
rect 574327 402972 574339 402984
rect 573524 402966 574339 402972
rect 573524 402965 574122 402966
rect 560128 402714 560134 402872
rect 560270 402714 560276 402872
rect 560128 402606 560276 402714
rect 566654 402747 575040 402867
rect 560128 402458 560726 402606
rect 566654 402584 566774 402747
rect 565664 402464 566774 402584
rect 565750 360473 573810 360593
rect 565750 358902 565870 360473
rect 566284 359987 566508 360011
rect 566278 359981 566524 359987
rect 566278 359801 566311 359981
rect 566491 359801 566524 359981
rect 566278 359795 566524 359801
rect 566284 359646 566508 359795
rect 559716 358047 560116 358061
rect 559716 357867 559740 358047
rect 559920 357867 560116 358047
rect 559716 357853 560116 357867
rect 559746 357568 559942 357853
rect 566292 357584 566447 359646
rect 573602 359359 573810 360473
rect 580266 359915 580370 359943
rect 580256 359913 580382 359915
rect 580256 359861 580293 359913
rect 580345 359861 580382 359913
rect 580256 359849 580382 359861
rect 580256 359797 580293 359849
rect 580345 359797 580382 359849
rect 580256 359795 580382 359797
rect 573602 359265 575010 359359
rect 573604 359239 575010 359265
rect 573604 357974 573842 359239
rect 573523 357968 573842 357974
rect 573523 357920 573925 357968
rect 573523 357612 573569 357920
rect 573877 357819 573925 357920
rect 580266 357926 580370 359795
rect 580266 357900 580464 357926
rect 573877 357818 574330 357819
rect 573877 357806 574338 357818
rect 573877 357612 574116 357806
rect 559732 357549 559942 357568
rect 566286 357578 566456 357584
rect 559732 357548 560116 357549
rect 559732 357542 560198 357548
rect 559732 357429 560070 357542
rect 559732 357122 559852 357429
rect 560058 357426 560070 357429
rect 560186 357426 560198 357542
rect 566286 357438 566298 357578
rect 566444 357438 566456 357578
rect 573523 357573 574116 357612
rect 574110 357570 574116 357573
rect 574332 357570 574338 357806
rect 580266 357714 580280 357900
rect 580448 357714 580464 357900
rect 580266 357708 580464 357714
rect 580274 357702 580454 357708
rect 574110 357558 574338 357570
rect 566286 357432 566456 357438
rect 560058 357420 560198 357426
rect 574592 357239 574712 357406
rect 566716 357124 574712 357239
rect 559732 357002 560730 357122
rect 565792 357119 574712 357124
rect 565792 357004 566836 357119
rect 508600 356609 508756 356611
rect 508600 356429 508620 356609
rect 508736 356429 508756 356609
rect 508600 356427 508756 356429
rect 565612 314307 573784 314427
rect 565612 313036 565732 314307
rect 566130 313806 566370 313813
rect 566130 313680 566160 313806
rect 566128 313626 566160 313680
rect 566340 313803 566370 313806
rect 566340 313626 566376 313803
rect 559656 311739 560258 311753
rect 559656 311559 559680 311739
rect 559860 311726 560258 311739
rect 559860 311568 560056 311726
rect 560246 311568 560258 311726
rect 559860 311559 560258 311568
rect 559656 311557 560258 311559
rect 566128 311694 566376 313626
rect 573560 313191 573784 314307
rect 580858 313787 580962 313791
rect 580770 313779 580962 313787
rect 580762 313774 580968 313779
rect 580762 313753 581008 313774
rect 580762 313637 580775 313753
rect 580955 313637 581008 313753
rect 580762 313611 581008 313637
rect 580770 313366 581008 313611
rect 574642 313191 575272 313296
rect 573560 313176 575272 313191
rect 573560 313071 574762 313176
rect 573560 311751 573814 313071
rect 580782 311865 581008 313366
rect 580509 311816 581008 311865
rect 580509 311812 580536 311816
rect 566128 311558 566156 311694
rect 559656 311545 560092 311557
rect 559662 311241 559894 311545
rect 566144 311508 566156 311558
rect 566358 311558 566376 311694
rect 573446 311691 574060 311751
rect 566358 311508 566370 311558
rect 566144 311502 566370 311508
rect 573446 311447 573523 311691
rect 573831 311599 574060 311691
rect 580507 311610 580536 311812
rect 580786 311610 581008 311816
rect 573831 311574 574728 311599
rect 580507 311590 581008 311610
rect 573831 311447 574558 311574
rect 573446 311410 574558 311447
rect 574718 311410 574728 311574
rect 573446 311401 574728 311410
rect 573446 311391 574064 311401
rect 574552 311398 574724 311401
rect 559662 311061 560868 311241
rect 575026 311181 575212 311292
rect 565562 311172 575212 311181
rect 565562 311061 575146 311172
<< via1 >>
rect 423872 691084 424132 691338
rect 476078 691094 476352 691356
rect 458146 689552 458266 689692
rect 406474 689426 406576 689524
rect 418238 688270 418324 688362
rect 465158 688228 465252 688344
rect 470582 688236 470670 688336
rect 413262 688056 413364 688162
rect 424234 688104 424342 688202
rect 476550 688050 476688 688184
rect 412022 686420 412170 686552
rect 463990 686390 464154 686542
rect 437516 668808 437660 668962
rect 446356 668822 446500 668974
rect 566340 583578 566492 583690
rect 580132 583568 580222 583676
rect 559788 581318 560010 581528
rect 573628 581122 573910 581438
rect 566210 507940 566316 507952
rect 566210 507840 566212 507940
rect 566212 507840 566310 507940
rect 566310 507840 566316 507940
rect 566210 507830 566316 507840
rect 559794 507678 559918 507792
rect 573616 507620 573914 507912
rect 580388 507856 580498 507968
rect 566197 449725 566377 449905
rect 559807 447937 559987 448117
rect 580848 449749 581028 449929
rect 573555 447499 573863 447743
rect 566283 405286 566463 405466
rect 559755 403231 559935 403347
rect 580116 405330 580168 405382
rect 573573 403001 573881 403309
rect 566311 359801 566491 359981
rect 559740 357867 559920 358047
rect 580293 359861 580345 359913
rect 580293 359797 580345 359849
rect 573569 357612 573877 357920
rect 508620 356429 508736 356609
rect 566160 313626 566340 313806
rect 559680 311559 559860 311739
rect 580775 313637 580955 313753
rect 573523 311447 573831 311691
<< metal2 >>
rect 476078 691356 476352 691366
rect 423872 691338 424132 691348
rect 476078 691084 476352 691094
rect 423872 691074 424132 691084
rect 458146 689692 458266 689702
rect 458146 689542 458266 689552
rect 406474 689524 406576 689534
rect 406474 689416 406576 689426
rect 418230 688374 418332 688384
rect 418230 688254 418332 688264
rect 465158 688344 465252 688354
rect 465158 688218 465252 688228
rect 470582 688336 470670 688346
rect 470582 688226 470670 688236
rect 424234 688202 424342 688212
rect 413252 688170 413372 688180
rect 424234 688094 424342 688104
rect 476550 688184 476688 688194
rect 413252 688034 413372 688044
rect 476550 688040 476688 688050
rect 412022 686552 412170 686562
rect 412022 686410 412170 686420
rect 463990 686542 464154 686552
rect 463990 686380 464154 686390
rect 446356 668974 446500 668984
rect 437516 668962 437660 668972
rect 446356 668812 446500 668822
rect 437516 668798 437660 668808
rect 566340 583690 566492 583700
rect 566340 583568 566492 583578
rect 580132 583676 580222 583686
rect 580132 583558 580222 583568
rect 559788 581528 560010 581538
rect 559788 581308 560010 581318
rect 573628 581438 573910 581448
rect 573628 581112 573910 581122
rect 580388 507968 580498 507978
rect 566210 507956 566316 507962
rect 566204 507952 566316 507956
rect 566204 507946 566210 507952
rect 566204 507830 566210 507838
rect 566204 507828 566316 507830
rect 566210 507820 566316 507828
rect 573616 507912 573914 507922
rect 559794 507792 559918 507802
rect 559794 507668 559918 507678
rect 580388 507846 580498 507856
rect 573616 507610 573914 507620
rect 580846 449929 581030 449955
rect 566176 449905 566398 449917
rect 566176 449883 566197 449905
rect 566377 449883 566398 449905
rect 566176 449747 566179 449883
rect 566395 449747 566398 449883
rect 566176 449725 566197 449747
rect 566377 449725 566398 449747
rect 566176 449713 566398 449725
rect 580846 449749 580848 449929
rect 581028 449749 581030 449929
rect 580846 449723 581030 449749
rect 559792 448117 560002 448143
rect 559792 447937 559807 448117
rect 559987 447937 560002 448117
rect 559792 447911 560002 447937
rect 573554 447743 573864 447767
rect 573554 447499 573555 447743
rect 573863 447499 573864 447743
rect 573554 447475 573864 447499
rect 566270 405484 566476 405495
rect 566270 405466 566305 405484
rect 566441 405466 566476 405484
rect 566270 405286 566283 405466
rect 566463 405286 566476 405466
rect 580088 405384 580196 405421
rect 580088 405328 580114 405384
rect 580170 405328 580196 405384
rect 580088 405291 580196 405328
rect 566270 405268 566305 405286
rect 566441 405268 566476 405286
rect 566270 405257 566476 405268
rect 559750 403357 559940 403387
rect 559750 403347 559777 403357
rect 559913 403347 559940 403357
rect 559750 403231 559755 403347
rect 559935 403231 559940 403347
rect 559750 403221 559777 403231
rect 559913 403221 559940 403231
rect 559750 403191 559940 403221
rect 573552 403309 573902 403331
rect 573552 403001 573573 403309
rect 573881 403001 573902 403309
rect 573552 402979 573902 403001
rect 541978 389509 542092 389529
rect 541978 389453 542007 389509
rect 542063 389453 542092 389509
rect 541978 389433 542092 389453
rect 541972 380673 542094 380687
rect 541972 380617 542005 380673
rect 542061 380617 542094 380673
rect 541972 380593 542094 380617
rect 541972 380537 542005 380593
rect 542061 380537 542094 380593
rect 541972 380523 542094 380537
rect 566288 359981 566514 359997
rect 566288 359959 566311 359981
rect 566491 359959 566514 359981
rect 566288 359823 566293 359959
rect 566509 359823 566514 359959
rect 566288 359801 566311 359823
rect 566491 359801 566514 359823
rect 566288 359785 566514 359801
rect 580266 359913 580372 359925
rect 580266 359883 580293 359913
rect 580345 359883 580372 359913
rect 580266 359827 580291 359883
rect 580347 359827 580372 359883
rect 580266 359797 580293 359827
rect 580345 359797 580372 359827
rect 580266 359785 580372 359797
rect 559726 358047 559934 358071
rect 559726 357867 559740 358047
rect 559920 357867 559934 358047
rect 559726 357843 559934 357867
rect 573554 357920 573892 357939
rect 573554 357612 573569 357920
rect 573877 357612 573892 357920
rect 573554 357593 573892 357612
rect 508610 356609 508746 356621
rect 508610 356587 508620 356609
rect 508736 356587 508746 356609
rect 508610 356429 508620 356451
rect 508736 356429 508746 356451
rect 508610 356417 508746 356429
rect 566140 313806 566360 313823
rect 566140 313784 566160 313806
rect 566340 313784 566360 313806
rect 566140 313648 566142 313784
rect 566358 313648 566360 313784
rect 566140 313626 566160 313648
rect 566340 313626 566360 313648
rect 566140 313609 566360 313626
rect 580772 313763 580958 313789
rect 580772 313753 580797 313763
rect 580933 313753 580958 313763
rect 580772 313637 580775 313753
rect 580955 313637 580958 313753
rect 580772 313627 580797 313637
rect 580933 313627 580958 313637
rect 580772 313601 580958 313627
rect 559666 311739 559874 311763
rect 559666 311559 559680 311739
rect 559860 311559 559874 311739
rect 559666 311535 559874 311559
rect 573506 311691 573848 311719
rect 573506 311447 573523 311691
rect 573831 311447 573848 311691
rect 573506 311419 573848 311447
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 423872 691084 424132 691338
rect 476078 691094 476352 691356
rect 458146 689552 458266 689692
rect 406474 689426 406576 689524
rect 418230 688362 418332 688374
rect 418230 688270 418238 688362
rect 418238 688270 418324 688362
rect 418324 688270 418332 688362
rect 418230 688264 418332 688270
rect 465158 688228 465252 688344
rect 470582 688236 470670 688336
rect 413252 688162 413372 688170
rect 413252 688056 413262 688162
rect 413262 688056 413364 688162
rect 413364 688056 413372 688162
rect 424234 688104 424342 688202
rect 413252 688044 413372 688056
rect 476550 688050 476688 688184
rect 412022 686420 412170 686552
rect 463990 686390 464154 686542
rect 437516 668808 437660 668962
rect 446356 668822 446500 668974
rect 566340 583578 566492 583690
rect 580132 583568 580222 583676
rect 559788 581318 560010 581528
rect 573628 581122 573910 581438
rect 566204 507838 566210 507946
rect 566210 507838 566316 507946
rect 559794 507678 559918 507792
rect 573616 507620 573914 507912
rect 580388 507856 580498 507968
rect 566179 449747 566197 449883
rect 566197 449747 566377 449883
rect 566377 449747 566395 449883
rect 580870 449771 581006 449907
rect 559829 447959 559965 448095
rect 573561 447513 573857 447729
rect 566305 405466 566441 405484
rect 566305 405286 566441 405466
rect 580114 405382 580170 405384
rect 580114 405330 580116 405382
rect 580116 405330 580168 405382
rect 580168 405330 580170 405382
rect 580114 405328 580170 405330
rect 566305 405268 566441 405286
rect 559777 403347 559913 403357
rect 559777 403231 559913 403347
rect 559777 403221 559913 403231
rect 573579 403007 573875 403303
rect 542007 389453 542063 389509
rect 542005 380617 542061 380673
rect 542005 380537 542061 380593
rect 566293 359823 566311 359959
rect 566311 359823 566491 359959
rect 566491 359823 566509 359959
rect 580291 359861 580293 359883
rect 580293 359861 580345 359883
rect 580345 359861 580347 359883
rect 580291 359849 580347 359861
rect 580291 359827 580293 359849
rect 580293 359827 580345 359849
rect 580345 359827 580347 359849
rect 559762 357889 559898 358025
rect 573575 357618 573871 357914
rect 508610 356451 508620 356587
rect 508620 356451 508736 356587
rect 508736 356451 508746 356587
rect 566142 313648 566160 313784
rect 566160 313648 566340 313784
rect 566340 313648 566358 313784
rect 580797 313753 580933 313763
rect 580797 313637 580933 313753
rect 580797 313627 580933 313637
rect 559702 311581 559838 311717
rect 573529 311461 573825 311677
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703482 418394 704800
rect 406344 691104 406354 691340
rect 406612 691104 406622 691340
rect 406404 689529 406584 691104
rect 406404 689524 406586 689529
rect 406404 689426 406474 689524
rect 406576 689426 406586 689524
rect 406404 689421 406586 689426
rect 406404 689412 406584 689421
rect 413128 688374 418426 703482
rect 465394 702876 470394 704800
rect 510594 703613 515394 704800
rect 423862 691338 424142 691343
rect 423862 691084 423872 691338
rect 424132 691084 424142 691338
rect 458040 691094 458050 691356
rect 458334 691094 458344 691356
rect 423862 691079 424142 691084
rect 458118 689692 458296 691094
rect 458118 689552 458146 689692
rect 458266 689552 458296 689692
rect 458118 689536 458296 689552
rect 413128 688264 418230 688374
rect 418332 688264 418426 688374
rect 413128 688170 418426 688264
rect 465042 688344 470794 702876
rect 510574 701285 515408 703613
rect 520594 703131 525394 704800
rect 510566 701189 515408 701285
rect 510566 700101 515400 701189
rect 520568 700588 525402 703131
rect 566594 702300 571594 704800
rect 510566 699600 515406 700101
rect 510550 698548 515406 699600
rect 520566 698548 525402 700588
rect 476068 691356 476362 691361
rect 476068 691094 476078 691356
rect 476352 691094 476362 691356
rect 476068 691089 476362 691094
rect 413128 688044 413252 688170
rect 413372 688044 418426 688170
rect 412012 686556 412180 686557
rect 412000 686414 412010 686556
rect 412174 686414 412184 686556
rect -800 680242 1700 685242
rect 413128 676163 418426 688044
rect 424190 688202 424390 688246
rect 424190 688104 424234 688202
rect 424342 688104 424390 688202
rect 424190 686560 424390 688104
rect 465042 688228 465158 688344
rect 465252 688336 470794 688344
rect 465252 688236 470582 688336
rect 470670 688236 470794 688336
rect 465252 688228 470794 688236
rect 424174 686342 424184 686560
rect 424398 686342 424408 686560
rect 463966 686368 463976 686548
rect 464170 686368 464180 686548
rect 413128 670865 438870 676163
rect 465042 676088 470794 688228
rect 476524 688184 476746 688212
rect 476524 688050 476550 688184
rect 476688 688050 476746 688184
rect 476524 686572 476746 688050
rect 510550 687360 515248 698548
rect 520566 687360 525388 698548
rect 510550 687048 515408 687360
rect 520566 687048 525404 687360
rect 476512 686390 476522 686572
rect 476744 686390 476754 686572
rect 510554 686489 515408 687048
rect 510554 686163 515388 686489
rect 510554 685661 510737 686163
rect 510576 678739 510737 685661
rect 515201 678739 515388 686163
rect 510576 678487 515388 678739
rect 520570 686139 525404 687048
rect 520570 678715 520737 686139
rect 525201 678715 525404 686139
rect 520570 678548 525404 678715
rect 582300 677984 584800 682984
rect 437480 668962 437708 670865
rect 445516 670336 470794 676088
rect 437480 668808 437516 668962
rect 437660 668808 437708 668962
rect 437480 668764 437708 668808
rect 446324 668974 446512 670336
rect 446324 668822 446356 668974
rect 446500 668822 446512 668974
rect 446324 668804 446512 668822
rect -800 643842 1660 648642
rect 567119 644605 581246 644615
rect 567119 644584 582932 644605
rect 567119 644323 584800 644584
rect 567119 640099 567336 644323
rect 573720 640099 584800 644323
rect 567119 639784 584800 640099
rect 567119 639769 582932 639784
rect -800 633842 1660 638642
rect 567322 634584 583190 634597
rect 567322 634265 584800 634584
rect 567310 634255 584800 634265
rect 567310 630031 567336 634255
rect 573720 630031 584800 634255
rect 567310 630021 584800 630031
rect 567322 629784 584800 630021
rect 567322 629761 583190 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 507976 583288 507986 583852
rect 508658 583674 508668 583852
rect 566330 583690 566502 583695
rect 566330 583674 566340 583690
rect 508658 583578 566340 583674
rect 566492 583674 566502 583690
rect 580122 583676 580232 583681
rect 580122 583674 580132 583676
rect 566492 583578 580132 583674
rect 508658 583568 580132 583578
rect 580222 583674 580232 583676
rect 580222 583568 584800 583674
rect 508658 583562 584800 583568
rect 508658 583288 508668 583562
rect 559778 581528 560020 581533
rect 559778 581318 559788 581528
rect 560010 581318 560020 581528
rect 559778 581313 560020 581318
rect 573618 581438 573920 581443
rect 573618 581122 573628 581438
rect 573910 581122 573920 581438
rect 573618 581117 573920 581122
rect 457252 565074 457262 571686
rect 463874 571176 574176 571686
rect 463874 565074 566918 571176
rect 458534 564368 566918 565074
rect 574066 564368 574176 571176
rect -800 559442 1660 564242
rect 458534 564226 574176 564368
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 552438 543310 552448 543448
rect 533090 536792 552448 543310
rect 559104 543310 559114 543448
rect 559104 536792 559862 543310
rect 582340 540562 584800 545362
rect 533090 536654 559862 536792
rect 457490 515352 457500 515868
rect -800 511530 480 511642
rect -800 510348 480 510460
rect 457142 509644 457500 515352
rect 463724 515352 463734 515868
rect 463724 509644 493426 515352
rect -800 509166 480 509278
rect -800 507984 480 508096
rect 457142 507742 493426 509644
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 457142 501632 457846 507742
rect 457836 501518 457846 501632
rect 464070 501632 493426 507742
rect 524200 513300 543128 513312
rect 524200 506708 554094 513300
rect 580380 507973 580582 507980
rect 580378 507968 580582 507973
rect 566200 507951 566210 507952
rect 566194 507946 566210 507951
rect 566194 507838 566204 507946
rect 566316 507944 566326 507952
rect 566194 507833 566210 507838
rect 566200 507830 566210 507833
rect 566316 507830 566412 507944
rect 559784 507792 559928 507797
rect 559784 507678 559794 507792
rect 559918 507678 559928 507792
rect 559784 507673 559928 507678
rect 566208 506708 566412 507830
rect 573606 507912 573924 507917
rect 573606 507620 573616 507912
rect 573914 507620 573924 507912
rect 580378 507856 580388 507968
rect 580498 507856 580582 507968
rect 580378 507851 580582 507856
rect 573606 507615 573924 507620
rect 580380 506708 580582 507851
rect 464070 501518 464080 501632
rect 524200 497912 581748 506708
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 544502 494257 581748 497912
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 544502 494252 583876 494257
rect 544502 494140 584800 494252
rect 544502 494133 583876 494140
rect 544502 492988 581748 494133
rect 533090 479346 553036 486002
rect 559692 479346 559702 486002
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect 457318 465204 457328 465550
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 456982 459326 457328 465204
rect 463552 465204 463562 465550
rect 463552 459326 567824 465204
rect 456982 458980 567824 459326
rect 574048 458980 574058 465204
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 566138 449883 566444 449929
rect 501842 449845 501966 449846
rect 566138 449845 566179 449883
rect 501842 449747 566179 449845
rect 566395 449845 566444 449883
rect 580836 449907 581040 449950
rect 580836 449845 580870 449907
rect 566395 449771 580870 449845
rect 581006 449845 581040 449907
rect 581006 449830 582616 449845
rect 581006 449771 584800 449830
rect 566395 449747 584800 449771
rect 501842 449721 584800 449747
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 501842 414997 501966 449721
rect 566138 449687 566444 449721
rect 582402 449718 584800 449721
rect 559782 448099 560012 448138
rect 559782 447955 559825 448099
rect 559969 447955 560012 448099
rect 559782 447916 560012 447955
rect 573544 447733 573874 447762
rect 573544 447509 573557 447733
rect 573861 447509 573874 447733
rect 573544 447480 573874 447509
rect 501016 414873 501966 414997
rect 501016 414809 501140 414873
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 566260 405484 566486 405490
rect 566260 405409 566305 405484
rect 542700 405297 566305 405409
rect 542700 389543 542812 405297
rect 566260 405268 566305 405297
rect 566441 405409 566486 405484
rect 580078 405409 580206 405416
rect 566441 405408 583886 405409
rect 566441 405384 584800 405408
rect 566441 405328 580114 405384
rect 580170 405328 584800 405384
rect 566441 405297 584800 405328
rect 566441 405268 566486 405297
rect 580078 405296 580206 405297
rect 583520 405296 584800 405297
rect 566260 405262 566486 405268
rect 559740 403361 559950 403382
rect 559740 403217 559773 403361
rect 559917 403217 559950 403361
rect 559740 403196 559950 403217
rect 573542 403307 573912 403326
rect 573542 403003 573575 403307
rect 573879 403003 573912 403307
rect 573542 402984 573912 403003
rect 541968 389509 542812 389543
rect 541968 389453 542007 389509
rect 542063 389453 542812 389509
rect 541968 389431 542812 389453
rect -800 381864 480 381976
rect -800 380682 480 380794
rect 541957 380673 545151 380712
rect 541957 380617 542005 380673
rect 542061 380624 545151 380673
rect 542061 380617 545155 380624
rect 541957 380593 545155 380617
rect 541957 380537 542005 380593
rect 542061 380537 545155 380593
rect 541957 380506 545155 380537
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 545037 359912 545155 380506
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 566278 359959 566524 359992
rect 566278 359912 566293 359959
rect 545037 359823 566293 359912
rect 566509 359912 566524 359959
rect 580256 359912 580382 359920
rect 566509 359883 580955 359912
rect 566509 359827 580291 359883
rect 580347 359827 580955 359883
rect 566509 359823 580955 359827
rect 545037 359794 580955 359823
rect 566278 359790 566524 359794
rect 580256 359790 580382 359794
rect 580837 358993 580955 359794
rect 580837 358986 583854 358993
rect 580837 358875 584800 358986
rect 580837 358868 580955 358875
rect 583520 358874 584800 358875
rect 559716 358029 559944 358066
rect 559716 357885 559758 358029
rect 559902 357885 559944 358029
rect 559716 357848 559944 357885
rect 573544 357918 573902 357934
rect 573544 357614 573571 357918
rect 573875 357614 573902 357918
rect 573544 357598 573902 357614
rect 508599 356587 509617 356620
rect 508599 356451 508610 356587
rect 508746 356451 509617 356587
rect 508599 356410 509617 356451
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 509407 313779 509617 356410
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 566130 313784 566370 313818
rect 566130 313779 566142 313784
rect 509407 313648 566142 313779
rect 566358 313779 566370 313784
rect 580762 313779 580968 313784
rect 566358 313764 583752 313779
rect 566358 313763 584800 313764
rect 566358 313648 580797 313763
rect 509407 313627 580797 313648
rect 580933 313652 584800 313763
rect 580933 313627 583887 313652
rect 509407 313602 583887 313627
rect 559656 311721 559884 311758
rect 559656 311577 559698 311721
rect 559842 311577 559884 311721
rect 559656 311540 559884 311577
rect 573496 311681 573858 311714
rect 573496 311457 573525 311681
rect 573829 311457 573858 311681
rect 573496 311424 573858 311457
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 406354 691104 406612 691340
rect 423872 691084 424132 691338
rect 458050 691094 458334 691356
rect 476078 691094 476352 691356
rect 412010 686552 412174 686556
rect 412010 686420 412022 686552
rect 412022 686420 412170 686552
rect 412170 686420 412174 686552
rect 412010 686414 412174 686420
rect 424184 686342 424398 686560
rect 463976 686542 464170 686548
rect 463976 686390 463990 686542
rect 463990 686390 464154 686542
rect 464154 686390 464170 686542
rect 463976 686368 464170 686390
rect 476522 686390 476744 686572
rect 510737 678739 515201 686163
rect 520737 678715 525201 686139
rect 567336 640099 573720 644323
rect 567336 630031 573720 634255
rect 507986 583288 508658 583852
rect 559788 581318 560010 581528
rect 573628 581122 573910 581438
rect 457262 565074 463874 571686
rect 566918 564368 574066 571176
rect 552448 536792 559104 543448
rect 457500 509644 463724 515868
rect 457846 501518 464070 507742
rect 566210 507946 566316 507952
rect 566210 507838 566316 507946
rect 566210 507830 566316 507838
rect 559794 507678 559918 507792
rect 573616 507620 573914 507912
rect 553036 479346 559692 486002
rect 457328 459326 463552 465550
rect 567824 458980 574048 465204
rect 559825 448095 559969 448099
rect 559825 447959 559829 448095
rect 559829 447959 559965 448095
rect 559965 447959 559969 448095
rect 559825 447955 559969 447959
rect 573557 447729 573861 447733
rect 573557 447513 573561 447729
rect 573561 447513 573857 447729
rect 573857 447513 573861 447729
rect 573557 447509 573861 447513
rect 559773 403357 559917 403361
rect 559773 403221 559777 403357
rect 559777 403221 559913 403357
rect 559913 403221 559917 403357
rect 559773 403217 559917 403221
rect 573575 403303 573879 403307
rect 573575 403007 573579 403303
rect 573579 403007 573875 403303
rect 573875 403007 573879 403303
rect 573575 403003 573879 403007
rect 559758 358025 559902 358029
rect 559758 357889 559762 358025
rect 559762 357889 559898 358025
rect 559898 357889 559902 358025
rect 559758 357885 559902 357889
rect 573571 357914 573875 357918
rect 573571 357618 573575 357914
rect 573575 357618 573871 357914
rect 573871 357618 573875 357914
rect 573571 357614 573875 357618
rect 559698 311717 559842 311721
rect 559698 311581 559702 311717
rect 559702 311581 559838 311717
rect 559838 311581 559842 311717
rect 559698 311577 559842 311581
rect 573525 311677 573829 311681
rect 573525 311461 573529 311677
rect 573529 311461 573825 311677
rect 573825 311461 573829 311677
rect 573525 311457 573829 311461
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 458049 691356 458335 691357
rect 406353 691340 406613 691341
rect 406353 691104 406354 691340
rect 406612 691104 406613 691340
rect 406353 691103 406613 691104
rect 424126 691338 424133 691339
rect 423871 691084 423872 691092
rect 424132 691084 424133 691338
rect 458049 691094 458050 691356
rect 458334 691094 458335 691356
rect 458049 691093 458335 691094
rect 476077 691356 476353 691357
rect 476077 691094 476078 691356
rect 476352 691094 476353 691356
rect 476077 691093 476353 691094
rect 423871 691083 424133 691084
rect 395910 686572 560048 686611
rect 395910 686560 476522 686572
rect 395910 686556 424184 686560
rect 395910 686414 412010 686556
rect 412174 686414 424184 686556
rect 395910 686342 424184 686414
rect 424398 686548 476522 686560
rect 424398 686368 463976 686548
rect 464170 686390 476522 686548
rect 476744 686390 560048 686572
rect 464170 686368 560048 686390
rect 424398 686342 560048 686368
rect 395910 686163 560048 686342
rect 395910 678739 510737 686163
rect 515201 686139 560048 686163
rect 515201 678739 520737 686139
rect 395910 678715 520737 678739
rect 525201 678715 560048 686139
rect 395910 678563 560048 678715
rect 406012 661332 407644 678563
rect 473960 662578 475592 678563
rect 406012 659700 414600 661332
rect 467972 660946 475592 662578
rect 507985 583852 508659 583853
rect 507985 583288 507986 583852
rect 508658 583288 508659 583852
rect 507985 583287 508659 583288
rect 457261 571686 463875 571687
rect 457261 565074 457262 571686
rect 463874 565074 463875 571686
rect 457261 565073 463875 565074
rect 457262 515868 463874 565073
rect 508046 547268 508622 583287
rect 551988 581528 560036 678563
rect 567319 644323 573737 644334
rect 567319 640099 567336 644323
rect 573720 640099 573737 644323
rect 567319 640088 573737 640099
rect 567319 634255 573737 634266
rect 567319 630031 567336 634255
rect 573720 630031 573737 634255
rect 567319 630020 573737 630031
rect 551988 581318 559788 581528
rect 560010 581318 560036 581528
rect 457262 509644 457500 515868
rect 463724 509644 463874 515868
rect 457262 507743 463874 509644
rect 551988 543448 560036 581318
rect 573627 581438 573911 581439
rect 573627 581122 573628 581438
rect 573910 581122 573911 581438
rect 573627 581121 573911 581122
rect 566917 571176 574067 571177
rect 566917 564368 566918 571176
rect 574066 564368 574067 571176
rect 566917 564367 574067 564368
rect 551988 536792 552448 543448
rect 559104 536792 560036 543448
rect 551988 507792 560036 536792
rect 566209 507952 566317 507953
rect 566209 507830 566210 507952
rect 566316 507830 566317 507952
rect 566209 507829 566317 507830
rect 573615 507912 573915 507913
rect 457262 507742 464071 507743
rect 457262 501518 457846 507742
rect 464070 501518 464071 507742
rect 457262 501517 464071 501518
rect 551988 507678 559794 507792
rect 559918 507678 560036 507792
rect 457262 465550 463874 501517
rect 457262 459996 457328 465550
rect 457327 459326 457328 459996
rect 463552 459996 463874 465550
rect 551988 486002 560036 507678
rect 573615 507620 573616 507912
rect 573914 507620 573915 507912
rect 573615 507619 573915 507620
rect 551988 479346 553036 486002
rect 559692 479346 560036 486002
rect 463552 459326 463553 459996
rect 457327 459325 463553 459326
rect 551988 451332 560036 479346
rect 567823 465204 574049 465205
rect 567823 458980 567824 465204
rect 574048 458980 574049 465204
rect 567823 458979 574049 458980
rect 551964 448099 560036 451332
rect 551964 447955 559825 448099
rect 559969 447955 560036 448099
rect 551964 444696 560036 447955
rect 573553 447739 573865 447758
rect 573553 447733 573591 447739
rect 573827 447733 573865 447739
rect 573553 447509 573557 447733
rect 573861 447509 573865 447733
rect 573553 447503 573591 447509
rect 573827 447503 573865 447509
rect 573553 447484 573865 447503
rect 551988 414063 560036 444696
rect 540426 412431 560036 414063
rect 551988 403361 560036 412431
rect 551988 403217 559773 403361
rect 559917 403217 560036 403361
rect 551988 359059 560036 403217
rect 573551 403307 573903 403322
rect 573551 403003 573575 403307
rect 573879 403003 573903 403307
rect 573551 402988 573903 403003
rect 534832 358029 560036 359059
rect 534832 357885 559758 358029
rect 559902 357885 560036 358029
rect 534832 357427 560036 357885
rect 573553 357918 573893 357930
rect 573553 357614 573571 357918
rect 573875 357614 573893 357918
rect 573553 357602 573893 357614
rect 551988 311721 560036 357427
rect 551988 311577 559698 311721
rect 559842 311577 560036 311721
rect 551988 154943 560036 311577
rect 573505 311687 573849 311710
rect 573505 311681 573559 311687
rect 573795 311681 573849 311687
rect 573505 311457 573525 311681
rect 573829 311457 573849 311681
rect 573505 311451 573559 311457
rect 573795 311451 573849 311457
rect 573505 311428 573849 311451
<< via4 >>
rect 406354 691104 406612 691340
rect 423866 691338 424126 691346
rect 423866 691092 423872 691338
rect 423872 691092 424126 691338
rect 458050 691094 458334 691356
rect 476078 691094 476352 691356
rect 567370 640173 573686 644249
rect 567370 630105 573686 634181
rect 573628 581122 573910 581438
rect 566918 564368 574066 571176
rect 573616 507620 573914 507912
rect 567824 458980 574048 465204
rect 573591 447733 573827 447739
rect 573591 447509 573827 447733
rect 573591 447503 573827 447509
rect 573609 403037 573845 403273
rect 573605 357648 573841 357884
rect 573559 311681 573795 311687
rect 573559 311457 573795 311681
rect 573559 311451 573795 311457
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 395311 691356 573934 697819
rect 395311 691346 458050 691356
rect 395311 691340 423866 691346
rect 395311 691104 406354 691340
rect 406612 691104 423866 691340
rect 395311 691092 423866 691104
rect 424126 691094 458050 691346
rect 458334 691094 476078 691356
rect 476352 691094 573934 691356
rect 424126 691092 573934 691094
rect 395311 691057 573934 691092
rect 398610 665680 400242 691057
rect 482026 665680 483658 691057
rect 398610 664048 421200 665680
rect 461900 664048 483658 665680
rect 567172 644249 573934 691057
rect 567172 640173 567370 644249
rect 573686 640173 573934 644249
rect 567172 634181 573934 640173
rect 567172 630105 567370 634181
rect 573686 630105 573934 634181
rect 567172 627323 573934 630105
rect 567170 621961 573956 627323
rect 567172 581438 573934 621961
rect 567172 581122 573628 581438
rect 573910 581122 573934 581438
rect 567172 571200 573934 581122
rect 566894 571176 574090 571200
rect 566894 564368 566918 571176
rect 574066 564368 574090 571176
rect 566894 564344 574090 564368
rect 567172 507936 573934 564344
rect 567172 507912 573938 507936
rect 567172 507620 573616 507912
rect 573914 507620 573938 507912
rect 567172 507596 573938 507620
rect 567172 465228 573934 507596
rect 567172 465204 574072 465228
rect 567172 458980 567824 465204
rect 574048 458980 574072 465204
rect 567172 458956 574072 458980
rect 567172 451332 573934 458956
rect 567148 447739 573934 451332
rect 567148 447503 573591 447739
rect 573827 447503 573934 447739
rect 567148 444696 573934 447503
rect 488794 422983 490426 423451
rect 567172 422983 573934 444696
rect 488794 421351 573934 422983
rect 488794 411215 490426 421351
rect 536998 420977 573934 421351
rect 537178 413157 538810 420977
rect 567172 403273 573934 420977
rect 567172 403037 573609 403273
rect 573845 403037 573934 403273
rect 488794 348933 490426 358653
rect 537178 348933 538810 359491
rect 567172 357884 573934 403037
rect 567172 357648 573605 357884
rect 573841 357648 573934 357884
rect 567172 348933 573934 357648
rect 488682 347301 573934 348933
rect 567172 311687 573934 347301
rect 567172 311451 573559 311687
rect 573795 311451 573934 311687
rect 567172 147394 573934 311451
use bandgaptop_flat_io  bandgaptop_flat_io_0
timestamp 1655695277
transform 0 1 -129800 -1 0 972356
box 422960 603262 502000 669400
use bgr_final  bgr_final_0
timestamp 1655699098
transform 0 -1 542076 -1 0 414982
box 0 0 58512 56576
use bgr_gen_8  bgr_gen_8_0
timestamp 1655764969
transform 1 0 412068 0 -1 668944
box 0 0 58512 56576
use nmos_flat  nmos_flat_0
timestamp 1655700407
transform -1 0 563137 0 1 358066
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_1
timestamp 1655700407
transform -1 0 563071 0 1 312130
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_2
timestamp 1655700407
transform -1 0 563201 0 1 403534
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_3
timestamp 1655700407
transform -1 0 563167 0 1 448522
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_4
timestamp 1655700407
transform -1 0 563375 0 1 582166
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_5
timestamp 1655700407
transform -1 0 563303 0 1 508484
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_6
timestamp 1655700407
transform 1 0 421454 0 1 688918
box -2706 -1060 2635 940
use nmos_flat  nmos_flat_7
timestamp 1655700407
transform 1 0 473730 0 1 688884
box -2706 -1060 2635 940
use pmos_flat  pmos_flat_0
timestamp 1655503347
transform -1 0 577475 0 1 448328
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_1
timestamp 1655503347
transform -1 0 577193 0 1 403846
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_2
timestamp 1655503347
transform -1 0 577239 0 1 358420
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_3
timestamp 1655503347
transform -1 0 577669 0 1 312352
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_4
timestamp 1655503347
transform -1 0 577171 0 1 582062
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_5
timestamp 1655503347
transform -1 0 577403 0 1 508572
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_6
timestamp 1655503347
transform -1 0 409419 0 1 688768
box -2742 -1060 2645 940
use pmos_flat  pmos_flat_7
timestamp 1655503347
transform -1 0 461215 0 1 688930
box -2742 -1060 2645 940
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 41 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 42 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 43 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 44 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 45 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 46 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 47 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 48 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 49 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 50 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 51 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 52 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 53 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 54 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 55 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 56 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 57 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 58 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 59 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 60 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 61 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 62 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 63 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 64 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 65 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 66 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 67 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 68 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 69 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 70 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 71 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 72 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 73 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 74 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 75 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 76 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 77 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 78 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 79 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 80 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 81 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 85 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 86 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 87 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 88 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 89 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 90 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 91 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 92 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 93 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 94 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 95 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 96 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 97 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 98 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 99 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 100 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 101 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 102 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 103 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 104 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 105 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 106 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 107 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 108 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 109 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 110 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 111 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 112 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 113 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 114 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 115 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 116 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 117 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 118 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 119 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 120 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 121 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 122 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 123 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 124 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 125 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 126 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 127 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 128 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 129 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 130 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 131 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 132 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 133 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 134 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 135 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 136 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 137 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 138 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 139 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 140 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 141 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 142 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 143 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 144 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 145 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 146 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 147 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 148 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 149 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 150 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 151 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 152 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 153 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 154 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 155 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 156 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 157 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 158 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 159 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 160 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 161 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 162 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 163 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 164 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 165 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 166 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 167 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 168 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 169 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 170 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 171 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 172 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 173 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 174 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 175 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 176 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 177 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 178 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 179 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 180 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 181 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 182 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 183 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 184 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 185 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 186 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 187 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 188 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 189 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 190 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 191 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 192 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 193 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 194 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 195 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 196 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 197 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 198 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 199 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 200 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 201 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 202 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 203 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 204 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 205 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 206 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 207 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 208 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 209 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 210 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 211 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 212 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 213 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 214 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 215 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 216 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 217 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 218 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 219 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 220 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 221 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 222 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 223 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 224 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 225 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 226 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 227 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 228 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 229 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 230 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 231 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 232 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 233 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 234 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 235 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 236 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 237 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 238 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 239 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 240 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 241 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 242 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 243 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 244 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 245 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 246 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 247 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 248 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 249 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 250 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 251 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 252 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 253 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 254 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 255 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 256 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 257 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 258 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 259 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 260 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 261 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 262 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 263 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 264 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 265 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 266 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 267 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 268 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 269 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 270 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 271 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 272 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 273 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 274 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 275 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 276 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 277 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 278 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 279 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 280 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 281 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 282 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 283 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 284 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 285 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 286 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 287 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 288 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 289 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 290 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 291 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 292 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 293 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 294 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 295 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 296 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 297 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 298 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 299 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 300 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 301 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 302 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 303 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 304 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 305 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 306 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 307 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 308 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 309 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 310 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 311 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 312 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 313 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 314 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 315 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 316 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 317 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 318 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 319 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 320 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 321 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 322 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 323 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 324 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 325 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 326 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 327 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 328 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 329 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 330 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 331 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 332 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 333 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 334 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 335 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 336 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 337 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 338 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 339 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 340 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 341 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 342 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 343 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 344 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 345 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 346 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 347 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 348 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 349 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 350 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 351 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 352 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 353 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 354 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 355 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 356 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 357 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 358 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 359 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 360 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 361 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 362 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 363 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 364 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 365 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 366 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 367 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 368 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 369 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 370 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 371 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 372 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 373 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 374 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 375 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 376 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 377 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 378 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 379 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 380 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 381 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 382 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 383 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 384 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 385 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 386 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 387 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 388 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 389 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 390 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 391 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 392 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 393 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 394 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 395 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 396 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 397 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 398 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 399 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 400 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 401 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 402 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 403 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 404 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 405 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 406 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 407 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 408 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 409 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 410 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 411 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 412 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 413 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 414 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 415 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 416 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 417 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 418 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 419 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 420 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 421 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 422 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 423 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 424 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 425 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 426 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 427 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 428 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 429 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 430 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 431 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 432 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 433 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 434 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 435 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 436 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 437 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 438 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 439 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 440 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 441 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 442 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 443 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 444 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 445 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 446 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 447 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 448 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 449 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 450 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 451 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 452 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 453 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 454 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 455 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 456 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 457 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 458 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 459 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 460 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 461 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 462 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 463 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 464 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 465 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 466 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 467 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 468 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 469 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 470 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 471 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 472 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 473 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 474 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 475 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 476 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 477 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 478 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 479 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 480 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 481 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 482 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 483 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 484 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 485 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 486 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 487 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 488 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 489 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 490 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 491 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 492 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 493 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 494 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 495 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 496 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 497 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 498 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 499 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 500 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 501 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 502 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 503 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 504 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 505 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 506 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 507 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 508 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 509 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 510 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 511 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 512 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 513 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 514 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 515 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 516 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 517 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 518 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 519 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 520 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 521 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 522 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 523 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 524 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 525 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 526 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 527 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 528 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 529 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 530 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 531 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 532 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 533 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 534 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 535 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 536 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 537 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 538 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 539 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 540 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 541 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 542 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 543 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 544 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 545 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 546 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 547 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 548 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 549 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 550 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 551 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 552 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 553 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 554 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 555 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 556 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 557 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 558 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 559 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 560 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 561 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 562 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 563 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 564 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 565 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 566 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 567 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 568 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 569 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 570 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 571 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 572 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 573 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 574 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 575 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 576 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 577 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 578 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 579 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 580 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 581 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 582 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 583 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 584 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 585 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 586 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 587 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 588 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 589 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 590 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 590 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 591 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 591 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 593 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 593 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 594 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 594 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 594 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 594 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 595 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 595 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 596 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 596 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 597 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 597 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 598 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 599 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 600 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 601 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 602 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 603 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 604 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 605 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 606 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 607 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 608 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 609 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 610 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 611 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 612 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 613 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 614 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 615 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 616 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 617 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 618 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 619 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 620 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 621 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 622 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 623 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 624 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 625 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 626 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 627 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 628 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 629 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 630 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 631 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 632 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 633 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 634 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 635 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 636 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 637 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 638 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 639 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 640 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 641 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 642 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 643 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 644 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 645 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 646 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 647 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 648 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 649 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 650 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 651 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 652 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 653 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 654 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 655 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 656 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 657 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 658 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 659 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 660 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 661 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 662 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 663 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 664 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 665 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 666 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 667 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 668 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 669 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 670 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 671 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 672 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 673 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 674 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 675 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 676 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 677 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 678 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 679 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 680 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 681 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 682 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 683 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 684 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 685 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 686 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 687 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 688 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 689 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 690 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 691 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 692 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 693 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 694 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 695 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 696 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 697 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 698 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 699 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 700 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 701 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 702 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 703 nsew
<< end >>
