magic
tech sky130A
magscale 1 2
timestamp 1655509990
<< nwell >>
rect 452648 637188 470026 637190
rect 442848 628688 452376 632030
rect 452648 629290 470914 637188
rect 452648 629288 458568 629290
rect 459358 629288 464068 629290
rect 464858 629288 470914 629290
<< pmoslvt >>
rect 443686 629350 444086 631930
rect 444258 629350 444658 631930
rect 444830 629350 445230 631930
rect 445402 629350 445802 631930
rect 445974 629350 446374 631930
rect 446546 629350 446946 631930
rect 447118 629350 447518 631930
rect 447690 629350 448090 631930
rect 448262 629350 448662 631930
rect 448834 629350 449234 631930
rect 449406 629350 449806 631930
rect 449978 629350 450378 631930
rect 450550 629350 450950 631930
rect 451122 629350 451522 631930
rect 453494 629388 453894 637128
rect 453952 629388 454352 637128
rect 454410 629388 454810 637128
rect 454868 629388 455268 637128
rect 455326 629388 455726 637128
rect 455784 629388 456184 637128
rect 456242 629388 456642 637128
rect 456700 629388 457100 637128
rect 457158 629388 457558 637128
rect 457616 629388 458016 637128
rect 458074 629388 458474 637128
rect 459452 629388 459852 637128
rect 459910 629388 460310 637128
rect 460368 629388 460768 637128
rect 460826 629388 461226 637128
rect 461284 629388 461684 637128
rect 461742 629388 462142 637128
rect 462200 629388 462600 637128
rect 462658 629388 463058 637128
rect 463116 629388 463516 637128
rect 463574 629388 463974 637128
rect 464952 629388 465352 637128
rect 465410 629388 465810 637128
rect 465868 629388 466268 637128
rect 466326 629388 466726 637128
rect 466784 629388 467184 637128
rect 467242 629388 467642 637128
rect 467700 629388 468100 637128
rect 468158 629388 468558 637128
rect 468616 629388 469016 637128
rect 469074 629388 469474 637128
rect 469532 629388 469932 637128
<< nmoslvt >>
rect 445072 636094 450472 636494
rect 440482 632820 440882 633220
rect 440940 632820 441340 633220
rect 441398 632820 441798 633220
rect 441856 632820 442256 633220
rect 442314 632820 442714 633220
rect 442772 632820 443172 633220
rect 445412 632542 445812 634342
rect 445984 632542 446384 634342
rect 446556 632542 446956 634342
rect 447128 632542 447528 634342
rect 447700 632542 448100 634342
rect 448272 632542 448672 634342
rect 448844 632542 449244 634342
rect 449416 632542 449816 634342
<< ndiff >>
rect 445072 636540 450472 636552
rect 445072 636506 445084 636540
rect 450460 636506 450472 636540
rect 445072 636494 450472 636506
rect 445072 636082 450472 636094
rect 445072 636048 445084 636082
rect 450460 636048 450472 636082
rect 445072 636036 450472 636048
rect 440424 633208 440482 633220
rect 440424 632832 440436 633208
rect 440470 632832 440482 633208
rect 440424 632820 440482 632832
rect 440882 633208 440940 633220
rect 440882 632832 440894 633208
rect 440928 632832 440940 633208
rect 440882 632820 440940 632832
rect 441340 633208 441398 633220
rect 441340 632832 441352 633208
rect 441386 632832 441398 633208
rect 441340 632820 441398 632832
rect 441798 633208 441856 633220
rect 441798 632832 441810 633208
rect 441844 632832 441856 633208
rect 441798 632820 441856 632832
rect 442256 633208 442314 633220
rect 442256 632832 442268 633208
rect 442302 632832 442314 633208
rect 442256 632820 442314 632832
rect 442714 633208 442772 633220
rect 442714 632832 442726 633208
rect 442760 632832 442772 633208
rect 442714 632820 442772 632832
rect 443172 633208 443230 633220
rect 443172 632832 443184 633208
rect 443218 632832 443230 633208
rect 443172 632820 443230 632832
rect 445354 634330 445412 634342
rect 445354 632554 445366 634330
rect 445400 632554 445412 634330
rect 445354 632542 445412 632554
rect 445812 634330 445870 634342
rect 445812 632554 445824 634330
rect 445858 632554 445870 634330
rect 445812 632542 445870 632554
rect 445926 634330 445984 634342
rect 445926 632554 445938 634330
rect 445972 632554 445984 634330
rect 445926 632542 445984 632554
rect 446384 634330 446442 634342
rect 446384 632554 446396 634330
rect 446430 632554 446442 634330
rect 446384 632542 446442 632554
rect 446498 634330 446556 634342
rect 446498 632554 446510 634330
rect 446544 632554 446556 634330
rect 446498 632542 446556 632554
rect 446956 634330 447014 634342
rect 446956 632554 446968 634330
rect 447002 632554 447014 634330
rect 446956 632542 447014 632554
rect 447070 634330 447128 634342
rect 447070 632554 447082 634330
rect 447116 632554 447128 634330
rect 447070 632542 447128 632554
rect 447528 634330 447586 634342
rect 447528 632554 447540 634330
rect 447574 632554 447586 634330
rect 447528 632542 447586 632554
rect 447642 634330 447700 634342
rect 447642 632554 447654 634330
rect 447688 632554 447700 634330
rect 447642 632542 447700 632554
rect 448100 634330 448158 634342
rect 448100 632554 448112 634330
rect 448146 632554 448158 634330
rect 448100 632542 448158 632554
rect 448214 634330 448272 634342
rect 448214 632554 448226 634330
rect 448260 632554 448272 634330
rect 448214 632542 448272 632554
rect 448672 634330 448730 634342
rect 448672 632554 448684 634330
rect 448718 632554 448730 634330
rect 448672 632542 448730 632554
rect 448786 634330 448844 634342
rect 448786 632554 448798 634330
rect 448832 632554 448844 634330
rect 448786 632542 448844 632554
rect 449244 634330 449302 634342
rect 449244 632554 449256 634330
rect 449290 632554 449302 634330
rect 449244 632542 449302 632554
rect 449358 634330 449416 634342
rect 449358 632554 449370 634330
rect 449404 632554 449416 634330
rect 449358 632542 449416 632554
rect 449816 634330 449874 634342
rect 449816 632554 449828 634330
rect 449862 632554 449874 634330
rect 449816 632542 449874 632554
<< pdiff >>
rect 453436 637116 453494 637128
rect 443628 631918 443686 631930
rect 443628 629362 443640 631918
rect 443674 629362 443686 631918
rect 443628 629350 443686 629362
rect 444086 631918 444144 631930
rect 444086 629362 444098 631918
rect 444132 629362 444144 631918
rect 444086 629350 444144 629362
rect 444200 631918 444258 631930
rect 444200 629362 444212 631918
rect 444246 629362 444258 631918
rect 444200 629350 444258 629362
rect 444658 631918 444716 631930
rect 444658 629362 444670 631918
rect 444704 629362 444716 631918
rect 444658 629350 444716 629362
rect 444772 631918 444830 631930
rect 444772 629362 444784 631918
rect 444818 629362 444830 631918
rect 444772 629350 444830 629362
rect 445230 631918 445288 631930
rect 445230 629362 445242 631918
rect 445276 629362 445288 631918
rect 445230 629350 445288 629362
rect 445344 631918 445402 631930
rect 445344 629362 445356 631918
rect 445390 629362 445402 631918
rect 445344 629350 445402 629362
rect 445802 631918 445860 631930
rect 445802 629362 445814 631918
rect 445848 629362 445860 631918
rect 445802 629350 445860 629362
rect 445916 631918 445974 631930
rect 445916 629362 445928 631918
rect 445962 629362 445974 631918
rect 445916 629350 445974 629362
rect 446374 631918 446432 631930
rect 446374 629362 446386 631918
rect 446420 629362 446432 631918
rect 446374 629350 446432 629362
rect 446488 631918 446546 631930
rect 446488 629362 446500 631918
rect 446534 629362 446546 631918
rect 446488 629350 446546 629362
rect 446946 631918 447004 631930
rect 446946 629362 446958 631918
rect 446992 629362 447004 631918
rect 446946 629350 447004 629362
rect 447060 631918 447118 631930
rect 447060 629362 447072 631918
rect 447106 629362 447118 631918
rect 447060 629350 447118 629362
rect 447518 631918 447576 631930
rect 447518 629362 447530 631918
rect 447564 629362 447576 631918
rect 447518 629350 447576 629362
rect 447632 631918 447690 631930
rect 447632 629362 447644 631918
rect 447678 629362 447690 631918
rect 447632 629350 447690 629362
rect 448090 631918 448148 631930
rect 448090 629362 448102 631918
rect 448136 629362 448148 631918
rect 448090 629350 448148 629362
rect 448204 631918 448262 631930
rect 448204 629362 448216 631918
rect 448250 629362 448262 631918
rect 448204 629350 448262 629362
rect 448662 631918 448720 631930
rect 448662 629362 448674 631918
rect 448708 629362 448720 631918
rect 448662 629350 448720 629362
rect 448776 631918 448834 631930
rect 448776 629362 448788 631918
rect 448822 629362 448834 631918
rect 448776 629350 448834 629362
rect 449234 631918 449292 631930
rect 449234 629362 449246 631918
rect 449280 629362 449292 631918
rect 449234 629350 449292 629362
rect 449348 631918 449406 631930
rect 449348 629362 449360 631918
rect 449394 629362 449406 631918
rect 449348 629350 449406 629362
rect 449806 631918 449864 631930
rect 449806 629362 449818 631918
rect 449852 629362 449864 631918
rect 449806 629350 449864 629362
rect 449920 631918 449978 631930
rect 449920 629362 449932 631918
rect 449966 629362 449978 631918
rect 449920 629350 449978 629362
rect 450378 631918 450436 631930
rect 450378 629362 450390 631918
rect 450424 629362 450436 631918
rect 450378 629350 450436 629362
rect 450492 631918 450550 631930
rect 450492 629362 450504 631918
rect 450538 629362 450550 631918
rect 450492 629350 450550 629362
rect 450950 631918 451008 631930
rect 450950 629362 450962 631918
rect 450996 629362 451008 631918
rect 450950 629350 451008 629362
rect 451064 631918 451122 631930
rect 451064 629362 451076 631918
rect 451110 629362 451122 631918
rect 451064 629350 451122 629362
rect 451522 631918 451580 631930
rect 451522 629362 451534 631918
rect 451568 629362 451580 631918
rect 453436 629400 453448 637116
rect 453482 629400 453494 637116
rect 453436 629388 453494 629400
rect 453894 637116 453952 637128
rect 453894 629400 453906 637116
rect 453940 629400 453952 637116
rect 453894 629388 453952 629400
rect 454352 637116 454410 637128
rect 454352 629400 454364 637116
rect 454398 629400 454410 637116
rect 454352 629388 454410 629400
rect 454810 637116 454868 637128
rect 454810 629400 454822 637116
rect 454856 629400 454868 637116
rect 454810 629388 454868 629400
rect 455268 637116 455326 637128
rect 455268 629400 455280 637116
rect 455314 629400 455326 637116
rect 455268 629388 455326 629400
rect 455726 637116 455784 637128
rect 455726 629400 455738 637116
rect 455772 629400 455784 637116
rect 455726 629388 455784 629400
rect 456184 637116 456242 637128
rect 456184 629400 456196 637116
rect 456230 629400 456242 637116
rect 456184 629388 456242 629400
rect 456642 637116 456700 637128
rect 456642 629400 456654 637116
rect 456688 629400 456700 637116
rect 456642 629388 456700 629400
rect 457100 637116 457158 637128
rect 457100 629400 457112 637116
rect 457146 629400 457158 637116
rect 457100 629388 457158 629400
rect 457558 637116 457616 637128
rect 457558 629400 457570 637116
rect 457604 629400 457616 637116
rect 457558 629388 457616 629400
rect 458016 637116 458074 637128
rect 458016 629400 458028 637116
rect 458062 629400 458074 637116
rect 458016 629388 458074 629400
rect 458474 637116 458532 637128
rect 458474 629400 458486 637116
rect 458520 629400 458532 637116
rect 459394 637116 459452 637128
rect 458474 629388 458532 629400
rect 459394 629400 459406 637116
rect 459440 629400 459452 637116
rect 459394 629388 459452 629400
rect 459852 637116 459910 637128
rect 459852 629400 459864 637116
rect 459898 629400 459910 637116
rect 459852 629388 459910 629400
rect 460310 637116 460368 637128
rect 460310 629400 460322 637116
rect 460356 629400 460368 637116
rect 460310 629388 460368 629400
rect 460768 637116 460826 637128
rect 460768 629400 460780 637116
rect 460814 629400 460826 637116
rect 460768 629388 460826 629400
rect 461226 637116 461284 637128
rect 461226 629400 461238 637116
rect 461272 629400 461284 637116
rect 461226 629388 461284 629400
rect 461684 637116 461742 637128
rect 461684 629400 461696 637116
rect 461730 629400 461742 637116
rect 461684 629388 461742 629400
rect 462142 637116 462200 637128
rect 462142 629400 462154 637116
rect 462188 629400 462200 637116
rect 462142 629388 462200 629400
rect 462600 637116 462658 637128
rect 462600 629400 462612 637116
rect 462646 629400 462658 637116
rect 462600 629388 462658 629400
rect 463058 637116 463116 637128
rect 463058 629400 463070 637116
rect 463104 629400 463116 637116
rect 463058 629388 463116 629400
rect 463516 637116 463574 637128
rect 463516 629400 463528 637116
rect 463562 629400 463574 637116
rect 463516 629388 463574 629400
rect 463974 637116 464032 637128
rect 463974 629400 463986 637116
rect 464020 629400 464032 637116
rect 464894 637116 464952 637128
rect 463974 629388 464032 629400
rect 464894 629400 464906 637116
rect 464940 629400 464952 637116
rect 464894 629388 464952 629400
rect 465352 637116 465410 637128
rect 465352 629400 465364 637116
rect 465398 629400 465410 637116
rect 465352 629388 465410 629400
rect 465810 637116 465868 637128
rect 465810 629400 465822 637116
rect 465856 629400 465868 637116
rect 465810 629388 465868 629400
rect 466268 637116 466326 637128
rect 466268 629400 466280 637116
rect 466314 629400 466326 637116
rect 466268 629388 466326 629400
rect 466726 637116 466784 637128
rect 466726 629400 466738 637116
rect 466772 629400 466784 637116
rect 466726 629388 466784 629400
rect 467184 637116 467242 637128
rect 467184 629400 467196 637116
rect 467230 629400 467242 637116
rect 467184 629388 467242 629400
rect 467642 637116 467700 637128
rect 467642 629400 467654 637116
rect 467688 629400 467700 637116
rect 467642 629388 467700 629400
rect 468100 637116 468158 637128
rect 468100 629400 468112 637116
rect 468146 629400 468158 637116
rect 468100 629388 468158 629400
rect 468558 637116 468616 637128
rect 468558 629400 468570 637116
rect 468604 629400 468616 637116
rect 468558 629388 468616 629400
rect 469016 637116 469074 637128
rect 469016 629400 469028 637116
rect 469062 629400 469074 637116
rect 469016 629388 469074 629400
rect 469474 637116 469532 637128
rect 469474 629400 469486 637116
rect 469520 629400 469532 637116
rect 469474 629388 469532 629400
rect 469932 637116 469990 637128
rect 469932 629400 469944 637116
rect 469978 629400 469990 637116
rect 469932 629388 469990 629400
rect 451522 629350 451580 629362
<< ndiffc >>
rect 445084 636506 450460 636540
rect 445084 636048 450460 636082
rect 440436 632832 440470 633208
rect 440894 632832 440928 633208
rect 441352 632832 441386 633208
rect 441810 632832 441844 633208
rect 442268 632832 442302 633208
rect 442726 632832 442760 633208
rect 443184 632832 443218 633208
rect 445366 632554 445400 634330
rect 445824 632554 445858 634330
rect 445938 632554 445972 634330
rect 446396 632554 446430 634330
rect 446510 632554 446544 634330
rect 446968 632554 447002 634330
rect 447082 632554 447116 634330
rect 447540 632554 447574 634330
rect 447654 632554 447688 634330
rect 448112 632554 448146 634330
rect 448226 632554 448260 634330
rect 448684 632554 448718 634330
rect 448798 632554 448832 634330
rect 449256 632554 449290 634330
rect 449370 632554 449404 634330
rect 449828 632554 449862 634330
<< pdiffc >>
rect 443640 629362 443674 631918
rect 444098 629362 444132 631918
rect 444212 629362 444246 631918
rect 444670 629362 444704 631918
rect 444784 629362 444818 631918
rect 445242 629362 445276 631918
rect 445356 629362 445390 631918
rect 445814 629362 445848 631918
rect 445928 629362 445962 631918
rect 446386 629362 446420 631918
rect 446500 629362 446534 631918
rect 446958 629362 446992 631918
rect 447072 629362 447106 631918
rect 447530 629362 447564 631918
rect 447644 629362 447678 631918
rect 448102 629362 448136 631918
rect 448216 629362 448250 631918
rect 448674 629362 448708 631918
rect 448788 629362 448822 631918
rect 449246 629362 449280 631918
rect 449360 629362 449394 631918
rect 449818 629362 449852 631918
rect 449932 629362 449966 631918
rect 450390 629362 450424 631918
rect 450504 629362 450538 631918
rect 450962 629362 450996 631918
rect 451076 629362 451110 631918
rect 451534 629362 451568 631918
rect 453448 629400 453482 637116
rect 453906 629400 453940 637116
rect 454364 629400 454398 637116
rect 454822 629400 454856 637116
rect 455280 629400 455314 637116
rect 455738 629400 455772 637116
rect 456196 629400 456230 637116
rect 456654 629400 456688 637116
rect 457112 629400 457146 637116
rect 457570 629400 457604 637116
rect 458028 629400 458062 637116
rect 458486 629400 458520 637116
rect 459406 629400 459440 637116
rect 459864 629400 459898 637116
rect 460322 629400 460356 637116
rect 460780 629400 460814 637116
rect 461238 629400 461272 637116
rect 461696 629400 461730 637116
rect 462154 629400 462188 637116
rect 462612 629400 462646 637116
rect 463070 629400 463104 637116
rect 463528 629400 463562 637116
rect 463986 629400 464020 637116
rect 464906 629400 464940 637116
rect 465364 629400 465398 637116
rect 465822 629400 465856 637116
rect 466280 629400 466314 637116
rect 466738 629400 466772 637116
rect 467196 629400 467230 637116
rect 467654 629400 467688 637116
rect 468112 629400 468146 637116
rect 468570 629400 468604 637116
rect 469028 629400 469062 637116
rect 469486 629400 469520 637116
rect 469944 629400 469978 637116
<< psubdiff >>
rect 437844 654854 483204 654878
rect 437844 653854 437868 654854
rect 483180 653854 483204 654854
rect 437844 653830 483204 653854
rect 482132 652830 483180 652854
rect 437892 652806 438940 652830
rect 437892 628654 437916 652806
rect 438916 628654 438940 652806
rect 440708 652724 451940 652748
rect 440708 651958 440732 652724
rect 451916 651958 451940 652724
rect 440708 651934 451940 651958
rect 452468 649188 453086 649212
rect 452468 642884 452492 649188
rect 453062 642884 453086 649188
rect 455712 649188 456330 649212
rect 452468 642860 453086 642884
rect 455712 642884 455736 649188
rect 456306 642884 456330 649188
rect 460672 649188 461290 649212
rect 455712 642860 456330 642884
rect 460672 642884 460696 649188
rect 461266 642884 461290 649188
rect 460672 642860 461290 642884
rect 475360 649188 475978 649212
rect 475360 642884 475384 649188
rect 475954 642884 475978 649188
rect 475360 642860 475978 642884
rect 482132 639936 482156 652830
rect 444342 637070 450842 637094
rect 444342 636738 444366 637070
rect 450818 636738 450842 637070
rect 444342 636714 450842 636738
rect 444764 634330 444964 634430
rect 439916 633524 443736 633548
rect 439916 633448 441330 633524
rect 442322 633448 443736 633524
rect 439916 633424 443736 633448
rect 439920 633370 440368 633424
rect 439920 632794 439944 633370
rect 440344 632794 440368 633370
rect 443286 633370 443734 633424
rect 443286 632794 443310 633370
rect 443710 632794 443734 633370
rect 439920 632770 440368 632794
rect 443286 632770 443734 632794
rect 444764 632730 444814 634330
rect 444914 632730 444964 634330
rect 444764 632630 444964 632730
rect 450264 634330 450464 634430
rect 450264 632730 450314 634330
rect 450414 632730 450464 634330
rect 450264 632630 450464 632730
rect 481152 629632 482156 639936
rect 437892 628630 438940 628654
rect 437868 627630 481156 627654
rect 437868 626630 437892 627630
rect 481132 626630 481156 627630
rect 437868 626606 481156 626630
rect 482132 626606 482156 629632
rect 483156 626606 483180 652830
rect 482132 626582 483180 626606
<< nsubdiff >>
rect 452748 636790 453348 636990
rect 442948 631830 443148 631930
rect 442948 629488 442998 631830
rect 443098 629488 443148 631830
rect 442948 629388 443148 629488
rect 452076 631830 452276 631930
rect 452076 629488 452126 631830
rect 452226 629488 452276 631830
rect 452748 629790 452948 636790
rect 453148 629790 453348 636790
rect 452748 629590 453348 629790
rect 452076 629388 452276 629488
rect 458658 636790 459258 636990
rect 458658 629790 458858 636790
rect 459058 629790 459258 636790
rect 458658 629590 459258 629790
rect 464158 636790 464758 636990
rect 464158 629790 464358 636790
rect 464558 629790 464758 636790
rect 464158 629590 464758 629790
rect 470114 636788 470714 636988
rect 470114 629788 470314 636788
rect 470514 629788 470714 636788
rect 470114 629588 470714 629788
rect 446480 628984 449022 629034
rect 446480 628884 446580 628984
rect 448922 628884 449022 628984
rect 446480 628834 449022 628884
<< psubdiffcont >>
rect 437868 653854 483180 654854
rect 437916 628654 438916 652806
rect 440732 651958 451916 652724
rect 452492 642884 453062 649188
rect 455736 642884 456306 649188
rect 460696 642884 461266 649188
rect 475384 642884 475954 649188
rect 444366 636738 450818 637070
rect 441330 633448 442322 633524
rect 439944 632794 440344 633370
rect 443310 632794 443710 633370
rect 444814 632730 444914 634330
rect 450314 632730 450414 634330
rect 437892 626630 481132 627630
rect 482156 626606 483156 652830
<< nsubdiffcont >>
rect 442998 629488 443098 631830
rect 452126 629488 452226 631830
rect 452948 629790 453148 636790
rect 458858 629790 459058 636790
rect 464358 629790 464558 636790
rect 470314 629788 470514 636788
rect 446580 628884 448922 628984
<< poly >>
rect 453494 637128 453894 637154
rect 453952 637128 454352 637154
rect 454410 637128 454810 637154
rect 454868 637128 455268 637154
rect 455326 637128 455726 637154
rect 455784 637128 456184 637154
rect 456242 637128 456642 637154
rect 456700 637128 457100 637154
rect 457158 637128 457558 637154
rect 457616 637128 458016 637154
rect 458074 637128 458474 637154
rect 459452 637128 459852 637154
rect 459910 637128 460310 637154
rect 460368 637128 460768 637154
rect 460826 637128 461226 637154
rect 461284 637128 461684 637154
rect 461742 637128 462142 637154
rect 462200 637128 462600 637154
rect 462658 637128 463058 637154
rect 463116 637128 463516 637154
rect 463574 637128 463974 637154
rect 464952 637128 465352 637154
rect 465410 637128 465810 637154
rect 465868 637128 466268 637154
rect 466326 637128 466726 637154
rect 466784 637128 467184 637154
rect 467242 637128 467642 637154
rect 467700 637128 468100 637154
rect 468158 637128 468558 637154
rect 468616 637128 469016 637154
rect 469074 637128 469474 637154
rect 469532 637128 469932 637154
rect 444984 636478 445072 636494
rect 444984 636110 445000 636478
rect 445034 636110 445072 636478
rect 444984 636094 445072 636110
rect 450472 636094 450498 636494
rect 445412 634414 445812 634430
rect 445412 634380 445428 634414
rect 445796 634380 445812 634414
rect 445412 634342 445812 634380
rect 445984 634414 446384 634430
rect 445984 634380 446000 634414
rect 446368 634380 446384 634414
rect 445984 634342 446384 634380
rect 446556 634414 446956 634430
rect 446556 634380 446572 634414
rect 446940 634380 446956 634414
rect 446556 634342 446956 634380
rect 447128 634414 447528 634430
rect 447128 634380 447144 634414
rect 447512 634380 447528 634414
rect 447128 634342 447528 634380
rect 447700 634414 448100 634430
rect 447700 634380 447716 634414
rect 448084 634380 448100 634414
rect 447700 634342 448100 634380
rect 448272 634414 448672 634430
rect 448272 634380 448288 634414
rect 448656 634380 448672 634414
rect 448272 634342 448672 634380
rect 448844 634414 449244 634430
rect 448844 634380 448860 634414
rect 449228 634380 449244 634414
rect 448844 634342 449244 634380
rect 449416 634414 449816 634430
rect 449416 634380 449432 634414
rect 449800 634380 449816 634414
rect 449416 634342 449816 634380
rect 440482 633292 440882 633308
rect 440482 633258 440498 633292
rect 440866 633258 440882 633292
rect 440482 633220 440882 633258
rect 440940 633292 441340 633308
rect 440940 633258 440956 633292
rect 441324 633258 441340 633292
rect 440940 633220 441340 633258
rect 441398 633292 441798 633308
rect 441398 633258 441414 633292
rect 441782 633258 441798 633292
rect 441398 633220 441798 633258
rect 441856 633292 442256 633308
rect 441856 633258 441872 633292
rect 442240 633258 442256 633292
rect 441856 633220 442256 633258
rect 442314 633292 442714 633308
rect 442314 633258 442330 633292
rect 442698 633258 442714 633292
rect 442314 633220 442714 633258
rect 442772 633292 443172 633308
rect 442772 633258 442788 633292
rect 443156 633258 443172 633292
rect 442772 633220 443172 633258
rect 440482 632794 440882 632820
rect 440940 632794 441340 632820
rect 441398 632794 441798 632820
rect 441856 632794 442256 632820
rect 442314 632794 442714 632820
rect 442772 632794 443172 632820
rect 445412 632516 445812 632542
rect 445984 632516 446384 632542
rect 446556 632516 446956 632542
rect 447128 632516 447528 632542
rect 447700 632516 448100 632542
rect 448272 632516 448672 632542
rect 448844 632516 449244 632542
rect 449416 632516 449816 632542
rect 443686 632011 444086 632027
rect 443686 631977 443702 632011
rect 444070 631977 444086 632011
rect 443686 631930 444086 631977
rect 444258 632011 444658 632027
rect 444258 631977 444274 632011
rect 444642 631977 444658 632011
rect 444258 631930 444658 631977
rect 444830 632011 445230 632027
rect 444830 631977 444846 632011
rect 445214 631977 445230 632011
rect 444830 631930 445230 631977
rect 445402 632011 445802 632027
rect 445402 631977 445418 632011
rect 445786 631977 445802 632011
rect 445402 631930 445802 631977
rect 445974 632011 446374 632027
rect 445974 631977 445990 632011
rect 446358 631977 446374 632011
rect 445974 631930 446374 631977
rect 446546 632011 446946 632027
rect 446546 631977 446562 632011
rect 446930 631977 446946 632011
rect 446546 631930 446946 631977
rect 447118 632011 447518 632027
rect 447118 631977 447134 632011
rect 447502 631977 447518 632011
rect 447118 631930 447518 631977
rect 447690 632011 448090 632027
rect 447690 631977 447706 632011
rect 448074 631977 448090 632011
rect 447690 631930 448090 631977
rect 448262 632011 448662 632027
rect 448262 631977 448278 632011
rect 448646 631977 448662 632011
rect 448262 631930 448662 631977
rect 448834 632011 449234 632027
rect 448834 631977 448850 632011
rect 449218 631977 449234 632011
rect 448834 631930 449234 631977
rect 449406 632011 449806 632027
rect 449406 631977 449422 632011
rect 449790 631977 449806 632011
rect 449406 631930 449806 631977
rect 449978 632011 450378 632027
rect 449978 631977 449994 632011
rect 450362 631977 450378 632011
rect 449978 631930 450378 631977
rect 450550 632011 450950 632027
rect 450550 631977 450566 632011
rect 450934 631977 450950 632011
rect 450550 631930 450950 631977
rect 451122 632011 451522 632027
rect 451122 631977 451138 632011
rect 451506 631977 451522 632011
rect 451122 631930 451522 631977
rect 443686 629324 444086 629350
rect 444258 629324 444658 629350
rect 444830 629324 445230 629350
rect 445402 629324 445802 629350
rect 445974 629324 446374 629350
rect 446546 629324 446946 629350
rect 447118 629324 447518 629350
rect 447690 629324 448090 629350
rect 448262 629324 448662 629350
rect 448834 629324 449234 629350
rect 449406 629324 449806 629350
rect 449978 629324 450378 629350
rect 450550 629324 450950 629350
rect 451122 629324 451522 629350
rect 453494 629341 453894 629388
rect 453494 629307 453510 629341
rect 453878 629307 453894 629341
rect 453494 629291 453894 629307
rect 453952 629341 454352 629388
rect 453952 629307 453968 629341
rect 454336 629307 454352 629341
rect 453952 629291 454352 629307
rect 454410 629341 454810 629388
rect 454410 629307 454426 629341
rect 454794 629307 454810 629341
rect 454410 629291 454810 629307
rect 454868 629341 455268 629388
rect 454868 629307 454884 629341
rect 455252 629307 455268 629341
rect 454868 629291 455268 629307
rect 455326 629341 455726 629388
rect 455326 629307 455342 629341
rect 455710 629307 455726 629341
rect 455326 629291 455726 629307
rect 455784 629341 456184 629388
rect 455784 629307 455800 629341
rect 456168 629307 456184 629341
rect 455784 629291 456184 629307
rect 456242 629341 456642 629388
rect 456242 629307 456258 629341
rect 456626 629307 456642 629341
rect 456242 629291 456642 629307
rect 456700 629341 457100 629388
rect 456700 629307 456716 629341
rect 457084 629307 457100 629341
rect 456700 629291 457100 629307
rect 457158 629341 457558 629388
rect 457158 629307 457174 629341
rect 457542 629307 457558 629341
rect 457158 629291 457558 629307
rect 457616 629341 458016 629388
rect 457616 629307 457632 629341
rect 458000 629307 458016 629341
rect 457616 629291 458016 629307
rect 458074 629341 458474 629388
rect 458074 629307 458090 629341
rect 458458 629307 458474 629341
rect 458074 629291 458474 629307
rect 459452 629341 459852 629388
rect 459452 629307 459468 629341
rect 459836 629307 459852 629341
rect 459452 629291 459852 629307
rect 459910 629341 460310 629388
rect 459910 629307 459926 629341
rect 460294 629307 460310 629341
rect 459910 629291 460310 629307
rect 460368 629341 460768 629388
rect 460368 629307 460384 629341
rect 460752 629307 460768 629341
rect 460368 629291 460768 629307
rect 460826 629341 461226 629388
rect 460826 629307 460842 629341
rect 461210 629307 461226 629341
rect 460826 629291 461226 629307
rect 461284 629341 461684 629388
rect 461284 629307 461300 629341
rect 461668 629307 461684 629341
rect 461284 629291 461684 629307
rect 461742 629341 462142 629388
rect 461742 629307 461758 629341
rect 462126 629307 462142 629341
rect 461742 629291 462142 629307
rect 462200 629341 462600 629388
rect 462200 629307 462216 629341
rect 462584 629307 462600 629341
rect 462200 629291 462600 629307
rect 462658 629341 463058 629388
rect 462658 629307 462674 629341
rect 463042 629307 463058 629341
rect 462658 629291 463058 629307
rect 463116 629341 463516 629388
rect 463116 629307 463132 629341
rect 463500 629307 463516 629341
rect 463116 629291 463516 629307
rect 463574 629341 463974 629388
rect 463574 629307 463590 629341
rect 463958 629307 463974 629341
rect 463574 629291 463974 629307
rect 464952 629341 465352 629388
rect 464952 629307 464968 629341
rect 465336 629307 465352 629341
rect 464952 629291 465352 629307
rect 465410 629341 465810 629388
rect 465410 629307 465426 629341
rect 465794 629307 465810 629341
rect 465410 629291 465810 629307
rect 465868 629341 466268 629388
rect 465868 629307 465884 629341
rect 466252 629307 466268 629341
rect 465868 629291 466268 629307
rect 466326 629341 466726 629388
rect 466326 629307 466342 629341
rect 466710 629307 466726 629341
rect 466326 629291 466726 629307
rect 466784 629341 467184 629388
rect 466784 629307 466800 629341
rect 467168 629307 467184 629341
rect 466784 629291 467184 629307
rect 467242 629341 467642 629388
rect 467242 629307 467258 629341
rect 467626 629307 467642 629341
rect 467242 629291 467642 629307
rect 467700 629341 468100 629388
rect 467700 629307 467716 629341
rect 468084 629307 468100 629341
rect 467700 629291 468100 629307
rect 468158 629341 468558 629388
rect 468158 629307 468174 629341
rect 468542 629307 468558 629341
rect 468158 629291 468558 629307
rect 468616 629341 469016 629388
rect 468616 629307 468632 629341
rect 469000 629307 469016 629341
rect 468616 629291 469016 629307
rect 469074 629341 469474 629388
rect 469074 629307 469090 629341
rect 469458 629307 469474 629341
rect 469074 629291 469474 629307
rect 469532 629341 469932 629388
rect 469532 629307 469548 629341
rect 469916 629307 469932 629341
rect 469532 629291 469932 629307
<< polycont >>
rect 445000 636110 445034 636478
rect 445428 634380 445796 634414
rect 446000 634380 446368 634414
rect 446572 634380 446940 634414
rect 447144 634380 447512 634414
rect 447716 634380 448084 634414
rect 448288 634380 448656 634414
rect 448860 634380 449228 634414
rect 449432 634380 449800 634414
rect 440498 633258 440866 633292
rect 440956 633258 441324 633292
rect 441414 633258 441782 633292
rect 441872 633258 442240 633292
rect 442330 633258 442698 633292
rect 442788 633258 443156 633292
rect 443702 631977 444070 632011
rect 444274 631977 444642 632011
rect 444846 631977 445214 632011
rect 445418 631977 445786 632011
rect 445990 631977 446358 632011
rect 446562 631977 446930 632011
rect 447134 631977 447502 632011
rect 447706 631977 448074 632011
rect 448278 631977 448646 632011
rect 448850 631977 449218 632011
rect 449422 631977 449790 632011
rect 449994 631977 450362 632011
rect 450566 631977 450934 632011
rect 451138 631977 451506 632011
rect 453510 629307 453878 629341
rect 453968 629307 454336 629341
rect 454426 629307 454794 629341
rect 454884 629307 455252 629341
rect 455342 629307 455710 629341
rect 455800 629307 456168 629341
rect 456258 629307 456626 629341
rect 456716 629307 457084 629341
rect 457174 629307 457542 629341
rect 457632 629307 458000 629341
rect 458090 629307 458458 629341
rect 459468 629307 459836 629341
rect 459926 629307 460294 629341
rect 460384 629307 460752 629341
rect 460842 629307 461210 629341
rect 461300 629307 461668 629341
rect 461758 629307 462126 629341
rect 462216 629307 462584 629341
rect 462674 629307 463042 629341
rect 463132 629307 463500 629341
rect 463590 629307 463958 629341
rect 464968 629307 465336 629341
rect 465426 629307 465794 629341
rect 465884 629307 466252 629341
rect 466342 629307 466710 629341
rect 466800 629307 467168 629341
rect 467258 629307 467626 629341
rect 467716 629307 468084 629341
rect 468174 629307 468542 629341
rect 468632 629307 469000 629341
rect 469090 629307 469458 629341
rect 469548 629307 469916 629341
<< xpolycontact >>
rect 456588 649250 457158 649682
rect 453316 647864 453886 648296
rect 453316 644108 453886 644540
rect 454134 647864 454704 648296
rect 454134 644108 454704 644540
rect 454952 647864 455522 648296
rect 454952 644108 455522 644540
rect 456588 644518 457158 644950
rect 457406 649250 457976 649682
rect 457406 644518 457976 644950
rect 458224 649250 458794 649682
rect 458224 644518 458794 644950
rect 459042 649250 459612 649682
rect 459042 644518 459612 644950
rect 461496 649188 462066 649620
rect 461496 642452 462066 642884
rect 462314 649188 462884 649620
rect 462314 642452 462884 642884
rect 463132 649188 463702 649620
rect 463132 642452 463702 642884
rect 463950 649188 464520 649620
rect 463950 642452 464520 642884
rect 464768 649188 465338 649620
rect 464768 642452 465338 642884
rect 465586 649188 466156 649620
rect 465586 642452 466156 642884
rect 466404 649188 466974 649620
rect 466404 642452 466974 642884
rect 467222 649188 467792 649620
rect 467222 642452 467792 642884
rect 468040 649188 468610 649620
rect 468040 642452 468610 642884
rect 468858 649188 469428 649620
rect 468858 642452 469428 642884
rect 469676 649188 470246 649620
rect 469676 642452 470246 642884
rect 470494 649188 471064 649620
rect 470494 642452 471064 642884
rect 471312 649188 471882 649620
rect 471312 642452 471882 642884
rect 472130 649188 472700 649620
rect 472130 642452 472700 642884
rect 472948 649188 473518 649620
rect 472948 642452 473518 642884
rect 473766 649188 474336 649620
rect 473766 642452 474336 642884
rect 474584 649188 475154 649620
rect 474584 642452 475154 642884
<< xpolyres >>
rect 453316 644540 453886 647864
rect 454134 644540 454704 647864
rect 454952 644540 455522 647864
rect 456588 644950 457158 649250
rect 457406 644950 457976 649250
rect 458224 644950 458794 649250
rect 459042 644950 459612 649250
rect 461496 642884 462066 649188
rect 462314 642884 462884 649188
rect 463132 642884 463702 649188
rect 463950 642884 464520 649188
rect 464768 642884 465338 649188
rect 465586 642884 466156 649188
rect 466404 642884 466974 649188
rect 467222 642884 467792 649188
rect 468040 642884 468610 649188
rect 468858 642884 469428 649188
rect 469676 642884 470246 649188
rect 470494 642884 471064 649188
rect 471312 642884 471882 649188
rect 472130 642884 472700 649188
rect 472948 642884 473518 649188
rect 473766 642884 474336 649188
rect 474584 642884 475154 649188
<< locali >>
rect 437844 654870 438868 654878
rect 437844 654854 438920 654870
rect 439020 654854 439144 654870
rect 439244 654854 439368 654870
rect 439468 654854 439592 654870
rect 439692 654854 439816 654870
rect 439916 654854 440040 654870
rect 440140 654854 440264 654870
rect 440364 654854 440488 654870
rect 440588 654854 440712 654870
rect 440812 654854 440936 654870
rect 441036 654854 441160 654870
rect 441260 654854 441384 654870
rect 441484 654854 441608 654870
rect 441708 654854 441832 654870
rect 441932 654854 442056 654870
rect 442156 654854 442280 654870
rect 442380 654854 442504 654870
rect 442604 654854 442728 654870
rect 442828 654854 442952 654870
rect 443052 654854 443176 654870
rect 443276 654854 443400 654870
rect 443500 654854 443624 654870
rect 443724 654854 443848 654870
rect 443948 654854 444072 654870
rect 444172 654854 444296 654870
rect 444396 654854 444520 654870
rect 444620 654854 444744 654870
rect 444844 654854 444968 654870
rect 445068 654854 445192 654870
rect 445292 654854 445416 654870
rect 445516 654854 449390 654870
rect 449490 654854 449614 654870
rect 449714 654854 449838 654870
rect 449938 654854 450062 654870
rect 450162 654854 450286 654870
rect 450386 654854 450510 654870
rect 450610 654854 450734 654870
rect 450834 654854 450958 654870
rect 451058 654854 451182 654870
rect 451282 654854 451406 654870
rect 451506 654854 451630 654870
rect 451730 654854 451854 654870
rect 451954 654854 452078 654870
rect 452178 654854 452302 654870
rect 452402 654854 452526 654870
rect 452626 654854 452750 654870
rect 452850 654854 452974 654870
rect 453074 654854 453198 654870
rect 453298 654854 453422 654870
rect 453522 654854 453646 654870
rect 453746 654854 453870 654870
rect 453970 654854 454094 654870
rect 454194 654854 454318 654870
rect 454418 654854 454542 654870
rect 454642 654854 454766 654870
rect 454866 654854 454990 654870
rect 455090 654854 455214 654870
rect 455314 654854 455438 654870
rect 455538 654854 455662 654870
rect 455762 654854 455886 654870
rect 455986 654854 475660 654870
rect 475760 654854 475884 654870
rect 475984 654854 476108 654870
rect 476208 654854 476332 654870
rect 476432 654854 476556 654870
rect 476656 654854 476780 654870
rect 476880 654854 477004 654870
rect 477104 654854 477228 654870
rect 477328 654854 477452 654870
rect 477552 654854 477676 654870
rect 477776 654854 477900 654870
rect 478000 654854 478124 654870
rect 478224 654854 478348 654870
rect 478448 654854 478572 654870
rect 478672 654854 478796 654870
rect 478896 654854 479020 654870
rect 479120 654854 479244 654870
rect 479344 654854 479468 654870
rect 479568 654854 479692 654870
rect 479792 654854 479916 654870
rect 480016 654854 480140 654870
rect 480240 654854 480364 654870
rect 480464 654854 480588 654870
rect 480688 654854 480812 654870
rect 480912 654854 481036 654870
rect 481136 654854 481260 654870
rect 481360 654854 481484 654870
rect 481584 654854 481708 654870
rect 481808 654854 481932 654870
rect 482032 654854 482156 654870
rect 482256 654854 483204 654878
rect 437844 653854 437868 654854
rect 483180 653854 483204 654854
rect 437844 653838 483204 653854
rect 437844 652822 438868 653838
rect 482204 652846 483204 653838
rect 482140 652830 483204 652846
rect 437844 652806 438932 652822
rect 437844 650178 437916 652806
rect 437844 650078 437894 650178
rect 437844 649954 437916 650078
rect 437844 649854 437894 649954
rect 437844 649730 437916 649854
rect 437844 649630 437894 649730
rect 437844 649506 437916 649630
rect 437844 649406 437894 649506
rect 437844 649282 437916 649406
rect 437844 649182 437894 649282
rect 437844 649058 437916 649182
rect 437844 648958 437894 649058
rect 437844 648834 437916 648958
rect 437844 648734 437894 648834
rect 437844 648610 437916 648734
rect 437844 648510 437894 648610
rect 437844 648386 437916 648510
rect 437844 648286 437894 648386
rect 437844 648162 437916 648286
rect 437844 648062 437894 648162
rect 437844 647938 437916 648062
rect 437844 647838 437894 647938
rect 437844 647714 437916 647838
rect 437844 647614 437894 647714
rect 437844 647490 437916 647614
rect 437844 647390 437894 647490
rect 437844 647266 437916 647390
rect 437844 647166 437894 647266
rect 437844 647042 437916 647166
rect 437844 646942 437894 647042
rect 437844 646818 437916 646942
rect 437844 646718 437894 646818
rect 437844 646594 437916 646718
rect 437844 646494 437894 646594
rect 437844 646370 437916 646494
rect 437844 646270 437894 646370
rect 437844 646146 437916 646270
rect 437844 646046 437894 646146
rect 437844 645922 437916 646046
rect 437844 645822 437894 645922
rect 437844 645698 437916 645822
rect 437844 645598 437894 645698
rect 437844 645474 437916 645598
rect 437844 645374 437894 645474
rect 437844 645250 437916 645374
rect 437844 645150 437894 645250
rect 437844 645026 437916 645150
rect 437844 644926 437894 645026
rect 437844 644802 437916 644926
rect 437844 644702 437894 644802
rect 437844 644578 437916 644702
rect 437844 644478 437894 644578
rect 437844 644354 437916 644478
rect 437844 644254 437894 644354
rect 437844 644130 437916 644254
rect 437844 644030 437894 644130
rect 437844 643906 437916 644030
rect 437844 643806 437894 643906
rect 437844 643682 437916 643806
rect 437844 643582 437894 643682
rect 437844 636778 437916 643582
rect 437844 636678 437894 636778
rect 437844 636554 437916 636678
rect 437844 636454 437894 636554
rect 437844 636330 437916 636454
rect 437844 636230 437894 636330
rect 437844 636106 437916 636230
rect 437844 636006 437894 636106
rect 437844 635882 437916 636006
rect 437844 635782 437894 635882
rect 437844 635658 437916 635782
rect 437844 635558 437894 635658
rect 437844 635434 437916 635558
rect 437844 635334 437894 635434
rect 437844 635210 437916 635334
rect 437844 635110 437894 635210
rect 437844 634986 437916 635110
rect 437844 634886 437894 634986
rect 437844 634762 437916 634886
rect 437844 634662 437894 634762
rect 437844 634538 437916 634662
rect 437844 634438 437894 634538
rect 437844 634314 437916 634438
rect 437844 634214 437894 634314
rect 437844 634090 437916 634214
rect 437844 633990 437894 634090
rect 437844 633866 437916 633990
rect 437844 633766 437894 633866
rect 437844 633642 437916 633766
rect 437844 633542 437894 633642
rect 437844 633418 437916 633542
rect 437844 633318 437894 633418
rect 437844 633194 437916 633318
rect 437844 633094 437894 633194
rect 437844 632970 437916 633094
rect 437844 632870 437894 632970
rect 437844 632746 437916 632870
rect 437844 632646 437894 632746
rect 437844 632522 437916 632646
rect 437844 632422 437894 632522
rect 437844 632298 437916 632422
rect 437844 632198 437894 632298
rect 437844 632074 437916 632198
rect 437844 631974 437894 632074
rect 437844 631850 437916 631974
rect 437844 631750 437894 631850
rect 437844 631626 437916 631750
rect 437844 631526 437894 631626
rect 437844 631402 437916 631526
rect 437844 631302 437894 631402
rect 437844 631178 437916 631302
rect 437844 631078 437894 631178
rect 437844 630954 437916 631078
rect 437844 630854 437894 630954
rect 437844 630730 437916 630854
rect 437844 630630 437894 630730
rect 437844 630506 437916 630630
rect 437844 630406 437894 630506
rect 437844 630282 437916 630406
rect 437844 630182 437894 630282
rect 437844 628654 437916 630182
rect 438916 628654 438932 652806
rect 455714 649250 456588 649682
rect 459612 649620 462066 649682
rect 459612 649250 461496 649620
rect 455714 649204 456318 649250
rect 452476 649188 453078 649204
rect 452476 648296 452492 649188
rect 452466 647854 452492 648296
rect 452476 643794 452492 647854
rect 452472 643290 452492 643794
rect 452476 642884 452492 643290
rect 453062 648296 453078 649188
rect 455714 649188 456322 649204
rect 459042 649188 461496 649250
rect 475154 649188 475978 649620
rect 455714 648692 455736 649188
rect 455720 648296 455736 648692
rect 453062 647864 453316 648296
rect 453886 647864 454134 648296
rect 454704 647864 454952 648296
rect 455522 647864 455736 648296
rect 453062 647854 455736 647864
rect 453062 643794 453078 647854
rect 455720 644540 455736 647854
rect 456306 644946 456322 649188
rect 460680 644950 460696 649188
rect 455522 644108 455736 644540
rect 453316 643798 453886 644108
rect 455720 643798 455736 644108
rect 456306 644518 456588 644946
rect 457158 644518 457264 644950
rect 458926 644518 459042 644950
rect 459612 644518 460696 644950
rect 456306 644420 457264 644518
rect 458926 644420 460696 644518
rect 453316 643794 455736 643798
rect 453062 643290 455736 643794
rect 453062 642884 453078 643290
rect 452476 642868 453078 642884
rect 455720 642884 455736 643290
rect 456306 643798 456322 644420
rect 456306 643290 456332 643798
rect 456306 642884 456322 643290
rect 460680 642884 460696 644420
rect 461266 642884 461282 649188
rect 475368 642884 475384 649188
rect 475954 642884 475970 649188
rect 455720 642868 456322 642884
rect 460672 642452 461496 642884
rect 475154 642452 475978 642884
rect 475771 639863 476241 639876
rect 477059 639863 477529 639876
rect 478347 639863 478817 639876
rect 479635 639863 480105 639876
rect 474953 639841 481008 639863
rect 474718 639701 481158 639841
rect 474718 638811 474953 639701
rect 475771 638811 476241 639701
rect 477059 638811 477529 639701
rect 478347 638811 478817 639701
rect 479635 638811 480105 639701
rect 480923 638811 481158 639701
rect 474718 638413 481158 638811
rect 474718 637523 474953 638413
rect 475771 637523 476241 638413
rect 477059 637523 477529 638413
rect 478347 637523 478817 638413
rect 479635 637523 480105 638413
rect 480923 637523 481158 638413
rect 453448 637116 453482 637132
rect 444350 637076 450834 637086
rect 444350 636732 444360 637076
rect 450824 636732 450834 637076
rect 444350 636722 450834 636732
rect 452748 636790 453348 636990
rect 445068 636506 445084 636540
rect 450460 636506 450476 636540
rect 445000 636478 445034 636494
rect 445000 636094 445034 636110
rect 445068 636048 445084 636082
rect 450460 636048 450476 636082
rect 445412 634380 445428 634414
rect 445796 634380 445812 634414
rect 445984 634380 446000 634414
rect 446368 634380 446384 634414
rect 446556 634380 446572 634414
rect 446940 634380 446956 634414
rect 447128 634380 447144 634414
rect 447512 634380 447528 634414
rect 447700 634380 447716 634414
rect 448084 634380 448100 634414
rect 448272 634380 448288 634414
rect 448656 634380 448672 634414
rect 448844 634380 448860 634414
rect 449228 634380 449244 634414
rect 449416 634380 449432 634414
rect 449800 634380 449816 634414
rect 444798 634330 444930 634346
rect 441314 633524 442338 633540
rect 441314 633448 441330 633524
rect 442322 633448 442338 633524
rect 441314 633408 442338 633448
rect 439928 633370 440360 633386
rect 439928 632794 439944 633370
rect 440344 633292 440360 633370
rect 441314 633356 441342 633408
rect 441394 633356 442258 633408
rect 442310 633356 442338 633408
rect 441314 633344 442338 633356
rect 443294 633370 443726 633386
rect 443294 633292 443310 633370
rect 440344 633258 440498 633292
rect 440866 633258 440882 633292
rect 440940 633258 440956 633292
rect 441324 633258 441414 633292
rect 441782 633258 441872 633292
rect 442240 633258 442330 633292
rect 442698 633258 442714 633292
rect 442772 633258 442788 633292
rect 443156 633258 443310 633292
rect 440344 633208 440470 633258
rect 440344 632832 440436 633208
rect 440344 632816 440470 632832
rect 440894 633208 440928 633224
rect 440894 632816 440928 632832
rect 441352 633208 441386 633224
rect 441352 632816 441386 632832
rect 441810 633208 441844 633224
rect 441810 632816 441844 632832
rect 442268 633208 442302 633224
rect 442268 632816 442302 632832
rect 442726 633208 442760 633224
rect 442726 632816 442760 632832
rect 443184 633208 443310 633258
rect 443218 632832 443310 633208
rect 443184 632816 443310 632832
rect 440344 632794 440360 632816
rect 439928 632778 440360 632794
rect 443294 632794 443310 632816
rect 443710 632794 443726 633370
rect 443294 632778 443726 632794
rect 444798 632730 444814 634330
rect 444914 632730 444930 634330
rect 444798 632714 444930 632730
rect 445366 634330 445400 634346
rect 445366 632538 445400 632554
rect 445824 634330 445858 634346
rect 445824 632538 445858 632554
rect 445938 634330 445972 634346
rect 445938 632538 445972 632554
rect 446396 634330 446430 634346
rect 446396 632538 446430 632554
rect 446510 634330 446544 634346
rect 446510 632538 446544 632554
rect 446968 634330 447002 634346
rect 446968 632538 447002 632554
rect 447082 634330 447116 634346
rect 447082 632538 447116 632554
rect 447540 634330 447574 634346
rect 447540 632538 447574 632554
rect 447654 634330 447688 634346
rect 447654 632538 447688 632554
rect 448112 634330 448146 634346
rect 448112 632538 448146 632554
rect 448226 634330 448260 634346
rect 448226 632538 448260 632554
rect 448684 634330 448718 634346
rect 448684 632538 448718 632554
rect 448798 634330 448832 634346
rect 448798 632538 448832 632554
rect 449256 634330 449290 634346
rect 449256 632538 449290 632554
rect 449370 634330 449404 634346
rect 449370 632538 449404 632554
rect 449828 634330 449862 634346
rect 450298 634330 450430 634346
rect 450298 632730 450314 634330
rect 450414 632730 450430 634330
rect 450298 632714 450430 632730
rect 449828 632538 449862 632554
rect 443686 631977 443702 632011
rect 444070 631977 444086 632011
rect 444258 631977 444274 632011
rect 444642 631977 444658 632011
rect 444830 631977 444846 632011
rect 445214 631977 445230 632011
rect 445402 631977 445418 632011
rect 445786 631977 445802 632011
rect 445974 631977 445990 632011
rect 446358 631977 446374 632011
rect 446546 631977 446562 632011
rect 446930 631977 446946 632011
rect 447118 631977 447134 632011
rect 447502 631977 447518 632011
rect 447690 631977 447706 632011
rect 448074 631977 448090 632011
rect 448262 631977 448278 632011
rect 448646 631977 448662 632011
rect 448834 631977 448850 632011
rect 449218 631977 449234 632011
rect 449406 631977 449422 632011
rect 449790 631977 449806 632011
rect 449978 631977 449994 632011
rect 450362 631977 450378 632011
rect 450550 631977 450566 632011
rect 450934 631977 450950 632011
rect 451122 631977 451138 632011
rect 451506 631977 451522 632011
rect 443640 631918 443674 631934
rect 442982 631830 443114 631842
rect 442982 629488 442998 631830
rect 443098 629488 443114 631830
rect 442982 629472 443114 629488
rect 443640 629346 443674 629362
rect 444098 631918 444132 631934
rect 444098 629346 444132 629362
rect 444212 631918 444246 631934
rect 444212 629346 444246 629362
rect 444670 631918 444704 631934
rect 444670 629346 444704 629362
rect 444784 631918 444818 631934
rect 444784 629346 444818 629362
rect 445242 631918 445276 631934
rect 445242 629346 445276 629362
rect 445356 631918 445390 631934
rect 445356 629346 445390 629362
rect 445814 631918 445848 631934
rect 445814 629346 445848 629362
rect 445928 631918 445962 631934
rect 445928 629346 445962 629362
rect 446386 631918 446420 631934
rect 446386 629346 446420 629362
rect 446500 631918 446534 631934
rect 446500 629346 446534 629362
rect 446958 631918 446992 631934
rect 446958 629346 446992 629362
rect 447072 631918 447106 631934
rect 447072 629346 447106 629362
rect 447530 631918 447564 631934
rect 447530 629346 447564 629362
rect 447644 631918 447678 631934
rect 447644 629346 447678 629362
rect 448102 631918 448136 631934
rect 448102 629346 448136 629362
rect 448216 631918 448250 631934
rect 448216 629346 448250 629362
rect 448674 631918 448708 631934
rect 448674 629346 448708 629362
rect 448788 631918 448822 631934
rect 448788 629346 448822 629362
rect 449246 631918 449280 631934
rect 449246 629346 449280 629362
rect 449360 631918 449394 631934
rect 449360 629346 449394 629362
rect 449818 631918 449852 631934
rect 449818 629346 449852 629362
rect 449932 631918 449966 631934
rect 449932 629346 449966 629362
rect 450390 631918 450424 631934
rect 450390 629346 450424 629362
rect 450504 631918 450538 631934
rect 450504 629346 450538 629362
rect 450962 631918 450996 631934
rect 450962 629346 450996 629362
rect 451076 631918 451110 631934
rect 451076 629346 451110 629362
rect 451534 631918 451568 631934
rect 452110 631830 452242 631842
rect 452110 629488 452126 631830
rect 452226 629488 452242 631830
rect 452110 629472 452242 629488
rect 452748 629790 452948 636790
rect 453148 629790 453348 636790
rect 451534 629346 451568 629362
rect 446568 628984 448938 629000
rect 446568 628884 446580 628984
rect 448922 628884 448938 628984
rect 446568 628868 448938 628884
rect 452748 628890 453348 629790
rect 453448 629384 453482 629400
rect 453906 637116 453940 637132
rect 453906 629384 453940 629400
rect 454364 637116 454398 637132
rect 454364 629384 454398 629400
rect 454822 637116 454856 637132
rect 454822 629384 454856 629400
rect 455280 637116 455314 637132
rect 455280 629384 455314 629400
rect 455738 637116 455772 637132
rect 455738 629384 455772 629400
rect 456196 637116 456230 637132
rect 456196 629384 456230 629400
rect 456654 637116 456688 637132
rect 456654 629384 456688 629400
rect 457112 637116 457146 637132
rect 457112 629384 457146 629400
rect 457570 637116 457604 637132
rect 457570 629384 457604 629400
rect 458028 637116 458062 637132
rect 458028 629384 458062 629400
rect 458486 637116 458520 637132
rect 459406 637116 459440 637132
rect 458486 629384 458520 629400
rect 458658 636790 459258 636990
rect 458658 629790 458858 636790
rect 459058 629790 459258 636790
rect 453494 629307 453510 629341
rect 453878 629307 453894 629341
rect 453952 629307 453968 629341
rect 454336 629307 454352 629341
rect 454410 629307 454426 629341
rect 454794 629307 454810 629341
rect 454868 629307 454884 629341
rect 455252 629307 455268 629341
rect 455326 629307 455342 629341
rect 455710 629307 455726 629341
rect 455784 629307 455800 629341
rect 456168 629307 456184 629341
rect 456242 629307 456258 629341
rect 456626 629307 456642 629341
rect 456700 629307 456716 629341
rect 457084 629307 457100 629341
rect 457158 629307 457174 629341
rect 457542 629307 457558 629341
rect 457616 629307 457632 629341
rect 458000 629307 458016 629341
rect 458074 629307 458090 629341
rect 458458 629307 458474 629341
rect 452748 628790 452848 628890
rect 453248 628790 453348 628890
rect 452748 628690 453348 628790
rect 458658 628890 459258 629790
rect 459406 629384 459440 629400
rect 459864 637116 459898 637132
rect 459864 629384 459898 629400
rect 460322 637116 460356 637132
rect 460322 629384 460356 629400
rect 460780 637116 460814 637132
rect 460780 629384 460814 629400
rect 461238 637116 461272 637132
rect 461238 629384 461272 629400
rect 461696 637116 461730 637132
rect 461696 629384 461730 629400
rect 462154 637116 462188 637132
rect 462154 629384 462188 629400
rect 462612 637116 462646 637132
rect 462612 629384 462646 629400
rect 463070 637116 463104 637132
rect 463070 629384 463104 629400
rect 463528 637116 463562 637132
rect 463528 629384 463562 629400
rect 463986 637116 464020 637132
rect 464906 637116 464940 637132
rect 463986 629384 464020 629400
rect 464158 636790 464758 636990
rect 464158 629790 464358 636790
rect 464558 629790 464758 636790
rect 459452 629307 459468 629341
rect 459836 629307 459852 629341
rect 459910 629307 459926 629341
rect 460294 629307 460310 629341
rect 460368 629307 460384 629341
rect 460752 629307 460768 629341
rect 460826 629307 460842 629341
rect 461210 629307 461226 629341
rect 461284 629307 461300 629341
rect 461668 629307 461684 629341
rect 461742 629307 461758 629341
rect 462126 629307 462142 629341
rect 462200 629307 462216 629341
rect 462584 629307 462600 629341
rect 462658 629307 462674 629341
rect 463042 629307 463058 629341
rect 463116 629307 463132 629341
rect 463500 629307 463516 629341
rect 463574 629307 463590 629341
rect 463958 629307 463974 629341
rect 458658 628790 458758 628890
rect 459158 628790 459258 628890
rect 458658 628690 459258 628790
rect 464158 628890 464758 629790
rect 464906 629384 464940 629400
rect 465364 637116 465398 637132
rect 465364 629384 465398 629400
rect 465822 637116 465856 637132
rect 465822 629384 465856 629400
rect 466280 637116 466314 637132
rect 466280 629384 466314 629400
rect 466738 637116 466772 637132
rect 466738 629384 466772 629400
rect 467196 637116 467230 637132
rect 467196 629384 467230 629400
rect 467654 637116 467688 637132
rect 467654 629384 467688 629400
rect 468112 637116 468146 637132
rect 468112 629384 468146 629400
rect 468570 637116 468604 637132
rect 468570 629384 468604 629400
rect 469028 637116 469062 637132
rect 469028 629384 469062 629400
rect 469486 637116 469520 637132
rect 469486 629384 469520 629400
rect 469944 637116 469978 637132
rect 474718 637125 481158 637523
rect 469944 629384 469978 629400
rect 470114 636788 470714 636988
rect 470114 629788 470314 636788
rect 470514 629788 470714 636788
rect 464952 629307 464968 629341
rect 465336 629307 465352 629341
rect 465410 629307 465426 629341
rect 465794 629307 465810 629341
rect 465868 629307 465884 629341
rect 466252 629307 466268 629341
rect 466326 629307 466342 629341
rect 466710 629307 466726 629341
rect 466784 629307 466800 629341
rect 467168 629307 467184 629341
rect 467242 629307 467258 629341
rect 467626 629307 467642 629341
rect 467700 629307 467716 629341
rect 468084 629307 468100 629341
rect 468158 629307 468174 629341
rect 468542 629307 468558 629341
rect 468616 629307 468632 629341
rect 469000 629307 469016 629341
rect 469074 629307 469090 629341
rect 469458 629307 469474 629341
rect 469532 629307 469548 629341
rect 469916 629307 469932 629341
rect 464158 628790 464258 628890
rect 464658 628790 464758 628890
rect 464158 628690 464758 628790
rect 470114 628888 470714 629788
rect 474718 636235 474953 637125
rect 475771 636235 476241 637125
rect 477059 636235 477529 637125
rect 478347 636235 478817 637125
rect 479635 636235 480105 637125
rect 480923 636235 481158 637125
rect 474718 635837 481158 636235
rect 474718 634947 474953 635837
rect 475771 634947 476241 635837
rect 477059 634947 477529 635837
rect 478347 634947 478817 635837
rect 479635 634947 480105 635837
rect 480923 634947 481158 635837
rect 474718 634549 481158 634947
rect 474718 633659 474953 634549
rect 475771 633659 476241 634549
rect 477059 633659 477529 634549
rect 478347 633659 478817 634549
rect 479635 633659 480105 634549
rect 480923 633659 481158 634549
rect 474718 633261 481158 633659
rect 474718 632371 474953 633261
rect 475771 632371 476241 633261
rect 477059 632371 477529 633261
rect 478347 632371 478817 633261
rect 479635 632371 480105 633261
rect 480923 632371 481158 633261
rect 474718 631973 481158 632371
rect 474718 631083 474953 631973
rect 475771 631083 476241 631973
rect 477059 631083 477529 631973
rect 478347 631083 478817 631973
rect 479635 631083 480105 631973
rect 480923 631083 481158 631973
rect 474718 630685 481158 631083
rect 474718 629867 474953 630685
rect 475771 629867 476241 630685
rect 477059 629867 477529 630685
rect 478347 629867 478817 630685
rect 479635 629867 480105 630685
rect 480923 629867 481158 630685
rect 474718 629731 481158 629867
rect 474718 629632 474953 629731
rect 475771 629632 476241 629731
rect 477059 629632 477529 629731
rect 478347 629632 478817 629731
rect 479635 629632 480105 629731
rect 480923 629632 481158 629731
rect 470114 628788 470214 628888
rect 470614 628788 470714 628888
rect 470114 628688 470714 628788
rect 437844 628638 438932 628654
rect 437844 627646 438868 628638
rect 437844 627630 438920 627646
rect 439020 627630 439144 627646
rect 439244 627630 439368 627646
rect 439468 627630 439592 627646
rect 439692 627630 439816 627646
rect 439916 627630 440040 627646
rect 440140 627630 440264 627646
rect 440364 627630 440488 627646
rect 440588 627630 440712 627646
rect 440812 627630 440936 627646
rect 441036 627630 441160 627646
rect 441260 627630 441384 627646
rect 441484 627630 441608 627646
rect 441708 627630 441832 627646
rect 441932 627630 442056 627646
rect 442156 627630 442280 627646
rect 442380 627630 442504 627646
rect 442604 627630 442728 627646
rect 442828 627630 442952 627646
rect 443052 627630 443176 627646
rect 443276 627630 443400 627646
rect 443500 627630 443624 627646
rect 443724 627630 443848 627646
rect 443948 627630 444072 627646
rect 444172 627630 444296 627646
rect 444396 627630 444520 627646
rect 444620 627630 444744 627646
rect 444844 627630 444968 627646
rect 445068 627630 445192 627646
rect 445292 627630 445416 627646
rect 445516 627630 449390 627646
rect 449490 627630 449614 627646
rect 449714 627630 449838 627646
rect 449938 627630 450062 627646
rect 450162 627630 450286 627646
rect 450386 627630 450510 627646
rect 450610 627630 450734 627646
rect 450834 627630 450958 627646
rect 451058 627630 451182 627646
rect 451282 627630 451406 627646
rect 451506 627630 451630 627646
rect 451730 627630 451854 627646
rect 451954 627630 452078 627646
rect 452178 627630 452302 627646
rect 452402 627630 452526 627646
rect 452626 627630 452750 627646
rect 452850 627630 452974 627646
rect 453074 627630 453198 627646
rect 453298 627630 453422 627646
rect 453522 627630 453646 627646
rect 453746 627630 453870 627646
rect 453970 627630 454094 627646
rect 454194 627630 454318 627646
rect 454418 627630 454542 627646
rect 454642 627630 454766 627646
rect 454866 627630 454990 627646
rect 455090 627630 455214 627646
rect 455314 627630 455438 627646
rect 455538 627630 455662 627646
rect 455762 627630 455886 627646
rect 455986 627630 475660 627646
rect 475760 627630 475884 627646
rect 475984 627630 476108 627646
rect 476208 627630 476332 627646
rect 476432 627630 476556 627646
rect 476656 627630 476780 627646
rect 476880 627630 477004 627646
rect 477104 627630 477228 627646
rect 477328 627630 477452 627646
rect 477552 627630 477676 627646
rect 477776 627630 477900 627646
rect 478000 627630 478124 627646
rect 478224 627630 478348 627646
rect 478448 627630 478572 627646
rect 478672 627630 478796 627646
rect 478896 627630 479020 627646
rect 479120 627630 479244 627646
rect 479344 627630 479468 627646
rect 479568 627630 479692 627646
rect 479792 627630 479916 627646
rect 480016 627630 480140 627646
rect 480240 627630 480364 627646
rect 480464 627630 480588 627646
rect 480688 627630 480812 627646
rect 480912 627630 481036 627646
rect 437844 626630 437892 627630
rect 481136 627606 481148 627646
rect 481136 627576 481260 627606
rect 481360 627576 481484 627606
rect 481584 627576 481708 627606
rect 481808 627576 481932 627606
rect 482140 627606 482156 652830
rect 483156 650178 483204 652830
rect 483170 650078 483204 650178
rect 483156 649954 483204 650078
rect 483170 649854 483204 649954
rect 483156 649730 483204 649854
rect 483170 649630 483204 649730
rect 483156 649506 483204 649630
rect 483170 649406 483204 649506
rect 483156 649282 483204 649406
rect 483170 649182 483204 649282
rect 483156 649058 483204 649182
rect 483170 648958 483204 649058
rect 483156 648834 483204 648958
rect 483170 648734 483204 648834
rect 483156 648610 483204 648734
rect 483170 648510 483204 648610
rect 483156 648386 483204 648510
rect 483170 648286 483204 648386
rect 483156 648162 483204 648286
rect 483170 648062 483204 648162
rect 483156 647938 483204 648062
rect 483170 647838 483204 647938
rect 483156 647714 483204 647838
rect 483170 647614 483204 647714
rect 483156 647490 483204 647614
rect 483170 647390 483204 647490
rect 483156 647266 483204 647390
rect 483170 647166 483204 647266
rect 483156 647042 483204 647166
rect 483170 646942 483204 647042
rect 483156 646818 483204 646942
rect 483170 646718 483204 646818
rect 483156 646594 483204 646718
rect 483170 646494 483204 646594
rect 483156 646370 483204 646494
rect 483170 646270 483204 646370
rect 483156 646146 483204 646270
rect 483170 646046 483204 646146
rect 483156 645922 483204 646046
rect 483170 645822 483204 645922
rect 483156 645698 483204 645822
rect 483170 645598 483204 645698
rect 483156 645474 483204 645598
rect 483170 645374 483204 645474
rect 483156 645250 483204 645374
rect 483170 645150 483204 645250
rect 483156 645026 483204 645150
rect 483170 644926 483204 645026
rect 483156 644802 483204 644926
rect 483170 644702 483204 644802
rect 483156 644578 483204 644702
rect 483170 644478 483204 644578
rect 483156 644354 483204 644478
rect 483170 644254 483204 644354
rect 483156 644130 483204 644254
rect 483170 644030 483204 644130
rect 483156 643906 483204 644030
rect 483170 643806 483204 643906
rect 483156 643682 483204 643806
rect 483170 643582 483204 643682
rect 483156 636778 483204 643582
rect 483170 636678 483204 636778
rect 483156 636554 483204 636678
rect 483170 636454 483204 636554
rect 483156 636330 483204 636454
rect 483170 636230 483204 636330
rect 483156 636106 483204 636230
rect 483170 636006 483204 636106
rect 483156 635882 483204 636006
rect 483170 635782 483204 635882
rect 483156 635658 483204 635782
rect 483170 635558 483204 635658
rect 483156 635434 483204 635558
rect 483170 635334 483204 635434
rect 483156 635210 483204 635334
rect 483170 635110 483204 635210
rect 483156 634986 483204 635110
rect 483170 634886 483204 634986
rect 483156 634762 483204 634886
rect 483170 634662 483204 634762
rect 483156 634538 483204 634662
rect 483170 634438 483204 634538
rect 483156 634314 483204 634438
rect 483170 634214 483204 634314
rect 483156 634090 483204 634214
rect 483170 633990 483204 634090
rect 483156 633866 483204 633990
rect 483170 633766 483204 633866
rect 483156 633642 483204 633766
rect 483170 633542 483204 633642
rect 483156 633418 483204 633542
rect 483170 633318 483204 633418
rect 483156 633194 483204 633318
rect 483170 633094 483204 633194
rect 483156 632970 483204 633094
rect 483170 632870 483204 632970
rect 483156 632746 483204 632870
rect 483170 632646 483204 632746
rect 483156 632522 483204 632646
rect 483170 632422 483204 632522
rect 483156 632298 483204 632422
rect 483170 632198 483204 632298
rect 483156 632074 483204 632198
rect 483170 631974 483204 632074
rect 483156 631850 483204 631974
rect 483170 631750 483204 631850
rect 483156 631626 483204 631750
rect 483170 631526 483204 631626
rect 483156 631402 483204 631526
rect 483170 631302 483204 631402
rect 483156 631178 483204 631302
rect 483170 631078 483204 631178
rect 483156 630954 483204 631078
rect 483170 630854 483204 630954
rect 483156 630730 483204 630854
rect 483170 630630 483204 630730
rect 483156 630506 483204 630630
rect 483170 630406 483204 630506
rect 483156 630282 483204 630406
rect 483170 630182 483204 630282
rect 482032 627576 482156 627606
rect 481132 627452 482156 627576
rect 481136 627352 481260 627452
rect 481360 627352 481484 627452
rect 481584 627352 481708 627452
rect 481808 627352 481932 627452
rect 482032 627352 482156 627452
rect 481132 627228 482156 627352
rect 481136 627128 481260 627228
rect 481360 627128 481484 627228
rect 481584 627128 481708 627228
rect 481808 627128 481932 627228
rect 482032 627128 482156 627228
rect 481132 627004 482156 627128
rect 481136 626904 481260 627004
rect 481360 626904 481484 627004
rect 481584 626904 481708 627004
rect 481808 626904 481932 627004
rect 482032 626904 482156 627004
rect 481132 626780 482156 626904
rect 481136 626680 481260 626780
rect 481360 626680 481484 626780
rect 481584 626680 481708 626780
rect 481808 626680 481932 626780
rect 482032 626680 482156 626780
rect 481132 626630 482156 626680
rect 437844 626614 482156 626630
rect 437844 626582 438868 626614
rect 480156 626606 482156 626614
rect 483156 626606 483204 630182
rect 480156 626582 483204 626606
<< viali >>
rect 438920 654854 439020 654876
rect 439144 654854 439244 654876
rect 439368 654854 439468 654876
rect 439592 654854 439692 654876
rect 439816 654854 439916 654876
rect 440040 654854 440140 654876
rect 440264 654854 440364 654876
rect 440488 654854 440588 654876
rect 440712 654854 440812 654876
rect 440936 654854 441036 654876
rect 441160 654854 441260 654876
rect 441384 654854 441484 654876
rect 441608 654854 441708 654876
rect 441832 654854 441932 654876
rect 442056 654854 442156 654876
rect 442280 654854 442380 654876
rect 442504 654854 442604 654876
rect 442728 654854 442828 654876
rect 442952 654854 443052 654876
rect 443176 654854 443276 654876
rect 443400 654854 443500 654876
rect 443624 654854 443724 654876
rect 443848 654854 443948 654876
rect 444072 654854 444172 654876
rect 444296 654854 444396 654876
rect 444520 654854 444620 654876
rect 444744 654854 444844 654876
rect 444968 654854 445068 654876
rect 445192 654854 445292 654876
rect 445416 654854 445516 654876
rect 449390 654854 449490 654876
rect 449614 654854 449714 654876
rect 449838 654854 449938 654876
rect 450062 654854 450162 654876
rect 450286 654854 450386 654876
rect 450510 654854 450610 654876
rect 450734 654854 450834 654876
rect 450958 654854 451058 654876
rect 451182 654854 451282 654876
rect 451406 654854 451506 654876
rect 451630 654854 451730 654876
rect 451854 654854 451954 654876
rect 452078 654854 452178 654876
rect 452302 654854 452402 654876
rect 452526 654854 452626 654876
rect 452750 654854 452850 654876
rect 452974 654854 453074 654876
rect 453198 654854 453298 654876
rect 453422 654854 453522 654876
rect 453646 654854 453746 654876
rect 453870 654854 453970 654876
rect 454094 654854 454194 654876
rect 454318 654854 454418 654876
rect 454542 654854 454642 654876
rect 454766 654854 454866 654876
rect 454990 654854 455090 654876
rect 455214 654854 455314 654876
rect 455438 654854 455538 654876
rect 455662 654854 455762 654876
rect 455886 654854 455986 654876
rect 475660 654854 475760 654896
rect 475884 654854 475984 654896
rect 476108 654854 476208 654896
rect 476332 654854 476432 654896
rect 476556 654854 476656 654896
rect 476780 654854 476880 654896
rect 477004 654854 477104 654896
rect 477228 654854 477328 654896
rect 477452 654854 477552 654896
rect 477676 654854 477776 654896
rect 477900 654854 478000 654896
rect 478124 654854 478224 654896
rect 478348 654854 478448 654896
rect 478572 654854 478672 654896
rect 478796 654854 478896 654896
rect 479020 654854 479120 654896
rect 479244 654854 479344 654896
rect 479468 654854 479568 654896
rect 479692 654854 479792 654896
rect 479916 654854 480016 654896
rect 480140 654854 480240 654896
rect 480364 654854 480464 654896
rect 480588 654854 480688 654896
rect 480812 654854 480912 654896
rect 481036 654854 481136 654896
rect 481260 654854 481360 654896
rect 481484 654854 481584 654896
rect 481708 654854 481808 654896
rect 481932 654854 482032 654896
rect 482156 654854 482256 654896
rect 438920 654776 439020 654854
rect 439144 654776 439244 654854
rect 439368 654776 439468 654854
rect 439592 654776 439692 654854
rect 439816 654776 439916 654854
rect 440040 654776 440140 654854
rect 440264 654776 440364 654854
rect 440488 654776 440588 654854
rect 440712 654776 440812 654854
rect 440936 654776 441036 654854
rect 441160 654776 441260 654854
rect 441384 654776 441484 654854
rect 441608 654776 441708 654854
rect 441832 654776 441932 654854
rect 442056 654776 442156 654854
rect 442280 654776 442380 654854
rect 442504 654776 442604 654854
rect 442728 654776 442828 654854
rect 442952 654776 443052 654854
rect 443176 654776 443276 654854
rect 443400 654776 443500 654854
rect 443624 654776 443724 654854
rect 443848 654776 443948 654854
rect 444072 654776 444172 654854
rect 444296 654776 444396 654854
rect 444520 654776 444620 654854
rect 444744 654776 444844 654854
rect 444968 654776 445068 654854
rect 445192 654776 445292 654854
rect 445416 654776 445516 654854
rect 449390 654776 449490 654854
rect 449614 654776 449714 654854
rect 449838 654776 449938 654854
rect 450062 654776 450162 654854
rect 450286 654776 450386 654854
rect 450510 654776 450610 654854
rect 450734 654776 450834 654854
rect 450958 654776 451058 654854
rect 451182 654776 451282 654854
rect 451406 654776 451506 654854
rect 451630 654776 451730 654854
rect 451854 654776 451954 654854
rect 452078 654776 452178 654854
rect 452302 654776 452402 654854
rect 452526 654776 452626 654854
rect 452750 654776 452850 654854
rect 452974 654776 453074 654854
rect 453198 654776 453298 654854
rect 453422 654776 453522 654854
rect 453646 654776 453746 654854
rect 453870 654776 453970 654854
rect 454094 654776 454194 654854
rect 454318 654776 454418 654854
rect 454542 654776 454642 654854
rect 454766 654776 454866 654854
rect 454990 654776 455090 654854
rect 455214 654776 455314 654854
rect 455438 654776 455538 654854
rect 455662 654776 455762 654854
rect 455886 654776 455986 654854
rect 475660 654796 475760 654854
rect 475884 654796 475984 654854
rect 476108 654796 476208 654854
rect 476332 654796 476432 654854
rect 476556 654796 476656 654854
rect 476780 654796 476880 654854
rect 477004 654796 477104 654854
rect 477228 654796 477328 654854
rect 477452 654796 477552 654854
rect 477676 654796 477776 654854
rect 477900 654796 478000 654854
rect 478124 654796 478224 654854
rect 478348 654796 478448 654854
rect 478572 654796 478672 654854
rect 478796 654796 478896 654854
rect 479020 654796 479120 654854
rect 479244 654796 479344 654854
rect 479468 654796 479568 654854
rect 479692 654796 479792 654854
rect 479916 654796 480016 654854
rect 480140 654796 480240 654854
rect 480364 654796 480464 654854
rect 480588 654796 480688 654854
rect 480812 654796 480912 654854
rect 481036 654796 481136 654854
rect 481260 654796 481360 654854
rect 481484 654796 481584 654854
rect 481708 654796 481808 654854
rect 481932 654796 482032 654854
rect 482156 654796 482256 654854
rect 438920 654552 439020 654652
rect 439144 654552 439244 654652
rect 439368 654552 439468 654652
rect 439592 654552 439692 654652
rect 439816 654552 439916 654652
rect 440040 654552 440140 654652
rect 440264 654552 440364 654652
rect 440488 654552 440588 654652
rect 440712 654552 440812 654652
rect 440936 654552 441036 654652
rect 441160 654552 441260 654652
rect 441384 654552 441484 654652
rect 441608 654552 441708 654652
rect 441832 654552 441932 654652
rect 442056 654552 442156 654652
rect 442280 654552 442380 654652
rect 442504 654552 442604 654652
rect 442728 654552 442828 654652
rect 442952 654552 443052 654652
rect 443176 654552 443276 654652
rect 443400 654552 443500 654652
rect 443624 654552 443724 654652
rect 443848 654552 443948 654652
rect 444072 654552 444172 654652
rect 444296 654552 444396 654652
rect 444520 654552 444620 654652
rect 444744 654552 444844 654652
rect 444968 654552 445068 654652
rect 445192 654552 445292 654652
rect 445416 654552 445516 654652
rect 449390 654552 449490 654652
rect 449614 654552 449714 654652
rect 449838 654552 449938 654652
rect 450062 654552 450162 654652
rect 450286 654552 450386 654652
rect 450510 654552 450610 654652
rect 450734 654552 450834 654652
rect 450958 654552 451058 654652
rect 451182 654552 451282 654652
rect 451406 654552 451506 654652
rect 451630 654552 451730 654652
rect 451854 654552 451954 654652
rect 452078 654552 452178 654652
rect 452302 654552 452402 654652
rect 452526 654552 452626 654652
rect 452750 654552 452850 654652
rect 452974 654552 453074 654652
rect 453198 654552 453298 654652
rect 453422 654552 453522 654652
rect 453646 654552 453746 654652
rect 453870 654552 453970 654652
rect 454094 654552 454194 654652
rect 454318 654552 454418 654652
rect 454542 654552 454642 654652
rect 454766 654552 454866 654652
rect 454990 654552 455090 654652
rect 455214 654552 455314 654652
rect 455438 654552 455538 654652
rect 455662 654552 455762 654652
rect 455886 654552 455986 654652
rect 475660 654572 475760 654672
rect 475884 654572 475984 654672
rect 476108 654572 476208 654672
rect 476332 654572 476432 654672
rect 476556 654572 476656 654672
rect 476780 654572 476880 654672
rect 477004 654572 477104 654672
rect 477228 654572 477328 654672
rect 477452 654572 477552 654672
rect 477676 654572 477776 654672
rect 477900 654572 478000 654672
rect 478124 654572 478224 654672
rect 478348 654572 478448 654672
rect 478572 654572 478672 654672
rect 478796 654572 478896 654672
rect 479020 654572 479120 654672
rect 479244 654572 479344 654672
rect 479468 654572 479568 654672
rect 479692 654572 479792 654672
rect 479916 654572 480016 654672
rect 480140 654572 480240 654672
rect 480364 654572 480464 654672
rect 480588 654572 480688 654672
rect 480812 654572 480912 654672
rect 481036 654572 481136 654672
rect 481260 654572 481360 654672
rect 481484 654572 481584 654672
rect 481708 654572 481808 654672
rect 481932 654572 482032 654672
rect 482156 654572 482256 654672
rect 438920 654328 439020 654428
rect 439144 654328 439244 654428
rect 439368 654328 439468 654428
rect 439592 654328 439692 654428
rect 439816 654328 439916 654428
rect 440040 654328 440140 654428
rect 440264 654328 440364 654428
rect 440488 654328 440588 654428
rect 440712 654328 440812 654428
rect 440936 654328 441036 654428
rect 441160 654328 441260 654428
rect 441384 654328 441484 654428
rect 441608 654328 441708 654428
rect 441832 654328 441932 654428
rect 442056 654328 442156 654428
rect 442280 654328 442380 654428
rect 442504 654328 442604 654428
rect 442728 654328 442828 654428
rect 442952 654328 443052 654428
rect 443176 654328 443276 654428
rect 443400 654328 443500 654428
rect 443624 654328 443724 654428
rect 443848 654328 443948 654428
rect 444072 654328 444172 654428
rect 444296 654328 444396 654428
rect 444520 654328 444620 654428
rect 444744 654328 444844 654428
rect 444968 654328 445068 654428
rect 445192 654328 445292 654428
rect 445416 654328 445516 654428
rect 449390 654328 449490 654428
rect 449614 654328 449714 654428
rect 449838 654328 449938 654428
rect 450062 654328 450162 654428
rect 450286 654328 450386 654428
rect 450510 654328 450610 654428
rect 450734 654328 450834 654428
rect 450958 654328 451058 654428
rect 451182 654328 451282 654428
rect 451406 654328 451506 654428
rect 451630 654328 451730 654428
rect 451854 654328 451954 654428
rect 452078 654328 452178 654428
rect 452302 654328 452402 654428
rect 452526 654328 452626 654428
rect 452750 654328 452850 654428
rect 452974 654328 453074 654428
rect 453198 654328 453298 654428
rect 453422 654328 453522 654428
rect 453646 654328 453746 654428
rect 453870 654328 453970 654428
rect 454094 654328 454194 654428
rect 454318 654328 454418 654428
rect 454542 654328 454642 654428
rect 454766 654328 454866 654428
rect 454990 654328 455090 654428
rect 455214 654328 455314 654428
rect 455438 654328 455538 654428
rect 455662 654328 455762 654428
rect 455886 654328 455986 654428
rect 475660 654348 475760 654448
rect 475884 654348 475984 654448
rect 476108 654348 476208 654448
rect 476332 654348 476432 654448
rect 476556 654348 476656 654448
rect 476780 654348 476880 654448
rect 477004 654348 477104 654448
rect 477228 654348 477328 654448
rect 477452 654348 477552 654448
rect 477676 654348 477776 654448
rect 477900 654348 478000 654448
rect 478124 654348 478224 654448
rect 478348 654348 478448 654448
rect 478572 654348 478672 654448
rect 478796 654348 478896 654448
rect 479020 654348 479120 654448
rect 479244 654348 479344 654448
rect 479468 654348 479568 654448
rect 479692 654348 479792 654448
rect 479916 654348 480016 654448
rect 480140 654348 480240 654448
rect 480364 654348 480464 654448
rect 480588 654348 480688 654448
rect 480812 654348 480912 654448
rect 481036 654348 481136 654448
rect 481260 654348 481360 654448
rect 481484 654348 481584 654448
rect 481708 654348 481808 654448
rect 481932 654348 482032 654448
rect 482156 654348 482256 654448
rect 438920 654104 439020 654204
rect 439144 654104 439244 654204
rect 439368 654104 439468 654204
rect 439592 654104 439692 654204
rect 439816 654104 439916 654204
rect 440040 654104 440140 654204
rect 440264 654104 440364 654204
rect 440488 654104 440588 654204
rect 440712 654104 440812 654204
rect 440936 654104 441036 654204
rect 441160 654104 441260 654204
rect 441384 654104 441484 654204
rect 441608 654104 441708 654204
rect 441832 654104 441932 654204
rect 442056 654104 442156 654204
rect 442280 654104 442380 654204
rect 442504 654104 442604 654204
rect 442728 654104 442828 654204
rect 442952 654104 443052 654204
rect 443176 654104 443276 654204
rect 443400 654104 443500 654204
rect 443624 654104 443724 654204
rect 443848 654104 443948 654204
rect 444072 654104 444172 654204
rect 444296 654104 444396 654204
rect 444520 654104 444620 654204
rect 444744 654104 444844 654204
rect 444968 654104 445068 654204
rect 445192 654104 445292 654204
rect 445416 654104 445516 654204
rect 449390 654104 449490 654204
rect 449614 654104 449714 654204
rect 449838 654104 449938 654204
rect 450062 654104 450162 654204
rect 450286 654104 450386 654204
rect 450510 654104 450610 654204
rect 450734 654104 450834 654204
rect 450958 654104 451058 654204
rect 451182 654104 451282 654204
rect 451406 654104 451506 654204
rect 451630 654104 451730 654204
rect 451854 654104 451954 654204
rect 452078 654104 452178 654204
rect 452302 654104 452402 654204
rect 452526 654104 452626 654204
rect 452750 654104 452850 654204
rect 452974 654104 453074 654204
rect 453198 654104 453298 654204
rect 453422 654104 453522 654204
rect 453646 654104 453746 654204
rect 453870 654104 453970 654204
rect 454094 654104 454194 654204
rect 454318 654104 454418 654204
rect 454542 654104 454642 654204
rect 454766 654104 454866 654204
rect 454990 654104 455090 654204
rect 455214 654104 455314 654204
rect 455438 654104 455538 654204
rect 455662 654104 455762 654204
rect 455886 654104 455986 654204
rect 475660 654124 475760 654224
rect 475884 654124 475984 654224
rect 476108 654124 476208 654224
rect 476332 654124 476432 654224
rect 476556 654124 476656 654224
rect 476780 654124 476880 654224
rect 477004 654124 477104 654224
rect 477228 654124 477328 654224
rect 477452 654124 477552 654224
rect 477676 654124 477776 654224
rect 477900 654124 478000 654224
rect 478124 654124 478224 654224
rect 478348 654124 478448 654224
rect 478572 654124 478672 654224
rect 478796 654124 478896 654224
rect 479020 654124 479120 654224
rect 479244 654124 479344 654224
rect 479468 654124 479568 654224
rect 479692 654124 479792 654224
rect 479916 654124 480016 654224
rect 480140 654124 480240 654224
rect 480364 654124 480464 654224
rect 480588 654124 480688 654224
rect 480812 654124 480912 654224
rect 481036 654124 481136 654224
rect 481260 654124 481360 654224
rect 481484 654124 481584 654224
rect 481708 654124 481808 654224
rect 481932 654124 482032 654224
rect 482156 654124 482256 654224
rect 438920 653880 439020 653980
rect 439144 653880 439244 653980
rect 439368 653880 439468 653980
rect 439592 653880 439692 653980
rect 439816 653880 439916 653980
rect 440040 653880 440140 653980
rect 440264 653880 440364 653980
rect 440488 653880 440588 653980
rect 440712 653880 440812 653980
rect 440936 653880 441036 653980
rect 441160 653880 441260 653980
rect 441384 653880 441484 653980
rect 441608 653880 441708 653980
rect 441832 653880 441932 653980
rect 442056 653880 442156 653980
rect 442280 653880 442380 653980
rect 442504 653880 442604 653980
rect 442728 653880 442828 653980
rect 442952 653880 443052 653980
rect 443176 653880 443276 653980
rect 443400 653880 443500 653980
rect 443624 653880 443724 653980
rect 443848 653880 443948 653980
rect 444072 653880 444172 653980
rect 444296 653880 444396 653980
rect 444520 653880 444620 653980
rect 444744 653880 444844 653980
rect 444968 653880 445068 653980
rect 445192 653880 445292 653980
rect 445416 653880 445516 653980
rect 449390 653880 449490 653980
rect 449614 653880 449714 653980
rect 449838 653880 449938 653980
rect 450062 653880 450162 653980
rect 450286 653880 450386 653980
rect 450510 653880 450610 653980
rect 450734 653880 450834 653980
rect 450958 653880 451058 653980
rect 451182 653880 451282 653980
rect 451406 653880 451506 653980
rect 451630 653880 451730 653980
rect 451854 653880 451954 653980
rect 452078 653880 452178 653980
rect 452302 653880 452402 653980
rect 452526 653880 452626 653980
rect 452750 653880 452850 653980
rect 452974 653880 453074 653980
rect 453198 653880 453298 653980
rect 453422 653880 453522 653980
rect 453646 653880 453746 653980
rect 453870 653880 453970 653980
rect 454094 653880 454194 653980
rect 454318 653880 454418 653980
rect 454542 653880 454642 653980
rect 454766 653880 454866 653980
rect 454990 653880 455090 653980
rect 455214 653880 455314 653980
rect 455438 653880 455538 653980
rect 455662 653880 455762 653980
rect 455886 653880 455986 653980
rect 475660 653900 475760 654000
rect 475884 653900 475984 654000
rect 476108 653900 476208 654000
rect 476332 653900 476432 654000
rect 476556 653900 476656 654000
rect 476780 653900 476880 654000
rect 477004 653900 477104 654000
rect 477228 653900 477328 654000
rect 477452 653900 477552 654000
rect 477676 653900 477776 654000
rect 477900 653900 478000 654000
rect 478124 653900 478224 654000
rect 478348 653900 478448 654000
rect 478572 653900 478672 654000
rect 478796 653900 478896 654000
rect 479020 653900 479120 654000
rect 479244 653900 479344 654000
rect 479468 653900 479568 654000
rect 479692 653900 479792 654000
rect 479916 653900 480016 654000
rect 480140 653900 480240 654000
rect 480364 653900 480464 654000
rect 480588 653900 480688 654000
rect 480812 653900 480912 654000
rect 481036 653900 481136 654000
rect 481260 653900 481360 654000
rect 481484 653900 481584 654000
rect 481708 653900 481808 654000
rect 481932 653900 482032 654000
rect 482156 653900 482256 654000
rect 437894 650078 437916 650178
rect 437916 650078 437994 650178
rect 438118 650078 438218 650178
rect 438342 650078 438442 650178
rect 438566 650078 438666 650178
rect 438790 650078 438890 650178
rect 437894 649854 437916 649954
rect 437916 649854 437994 649954
rect 438118 649854 438218 649954
rect 438342 649854 438442 649954
rect 438566 649854 438666 649954
rect 438790 649854 438890 649954
rect 437894 649630 437916 649730
rect 437916 649630 437994 649730
rect 438118 649630 438218 649730
rect 438342 649630 438442 649730
rect 438566 649630 438666 649730
rect 438790 649630 438890 649730
rect 437894 649406 437916 649506
rect 437916 649406 437994 649506
rect 438118 649406 438218 649506
rect 438342 649406 438442 649506
rect 438566 649406 438666 649506
rect 438790 649406 438890 649506
rect 437894 649182 437916 649282
rect 437916 649182 437994 649282
rect 438118 649182 438218 649282
rect 438342 649182 438442 649282
rect 438566 649182 438666 649282
rect 438790 649182 438890 649282
rect 437894 648958 437916 649058
rect 437916 648958 437994 649058
rect 438118 648958 438218 649058
rect 438342 648958 438442 649058
rect 438566 648958 438666 649058
rect 438790 648958 438890 649058
rect 437894 648734 437916 648834
rect 437916 648734 437994 648834
rect 438118 648734 438218 648834
rect 438342 648734 438442 648834
rect 438566 648734 438666 648834
rect 438790 648734 438890 648834
rect 437894 648510 437916 648610
rect 437916 648510 437994 648610
rect 438118 648510 438218 648610
rect 438342 648510 438442 648610
rect 438566 648510 438666 648610
rect 438790 648510 438890 648610
rect 437894 648286 437916 648386
rect 437916 648286 437994 648386
rect 438118 648286 438218 648386
rect 438342 648286 438442 648386
rect 438566 648286 438666 648386
rect 438790 648286 438890 648386
rect 437894 648062 437916 648162
rect 437916 648062 437994 648162
rect 438118 648062 438218 648162
rect 438342 648062 438442 648162
rect 438566 648062 438666 648162
rect 438790 648062 438890 648162
rect 437894 647838 437916 647938
rect 437916 647838 437994 647938
rect 438118 647838 438218 647938
rect 438342 647838 438442 647938
rect 438566 647838 438666 647938
rect 438790 647838 438890 647938
rect 437894 647614 437916 647714
rect 437916 647614 437994 647714
rect 438118 647614 438218 647714
rect 438342 647614 438442 647714
rect 438566 647614 438666 647714
rect 438790 647614 438890 647714
rect 437894 647390 437916 647490
rect 437916 647390 437994 647490
rect 438118 647390 438218 647490
rect 438342 647390 438442 647490
rect 438566 647390 438666 647490
rect 438790 647390 438890 647490
rect 437894 647166 437916 647266
rect 437916 647166 437994 647266
rect 438118 647166 438218 647266
rect 438342 647166 438442 647266
rect 438566 647166 438666 647266
rect 438790 647166 438890 647266
rect 437894 646942 437916 647042
rect 437916 646942 437994 647042
rect 438118 646942 438218 647042
rect 438342 646942 438442 647042
rect 438566 646942 438666 647042
rect 438790 646942 438890 647042
rect 437894 646718 437916 646818
rect 437916 646718 437994 646818
rect 438118 646718 438218 646818
rect 438342 646718 438442 646818
rect 438566 646718 438666 646818
rect 438790 646718 438890 646818
rect 437894 646494 437916 646594
rect 437916 646494 437994 646594
rect 438118 646494 438218 646594
rect 438342 646494 438442 646594
rect 438566 646494 438666 646594
rect 438790 646494 438890 646594
rect 437894 646270 437916 646370
rect 437916 646270 437994 646370
rect 438118 646270 438218 646370
rect 438342 646270 438442 646370
rect 438566 646270 438666 646370
rect 438790 646270 438890 646370
rect 437894 646046 437916 646146
rect 437916 646046 437994 646146
rect 438118 646046 438218 646146
rect 438342 646046 438442 646146
rect 438566 646046 438666 646146
rect 438790 646046 438890 646146
rect 437894 645822 437916 645922
rect 437916 645822 437994 645922
rect 438118 645822 438218 645922
rect 438342 645822 438442 645922
rect 438566 645822 438666 645922
rect 438790 645822 438890 645922
rect 437894 645598 437916 645698
rect 437916 645598 437994 645698
rect 438118 645598 438218 645698
rect 438342 645598 438442 645698
rect 438566 645598 438666 645698
rect 438790 645598 438890 645698
rect 437894 645374 437916 645474
rect 437916 645374 437994 645474
rect 438118 645374 438218 645474
rect 438342 645374 438442 645474
rect 438566 645374 438666 645474
rect 438790 645374 438890 645474
rect 437894 645150 437916 645250
rect 437916 645150 437994 645250
rect 438118 645150 438218 645250
rect 438342 645150 438442 645250
rect 438566 645150 438666 645250
rect 438790 645150 438890 645250
rect 437894 644926 437916 645026
rect 437916 644926 437994 645026
rect 438118 644926 438218 645026
rect 438342 644926 438442 645026
rect 438566 644926 438666 645026
rect 438790 644926 438890 645026
rect 437894 644702 437916 644802
rect 437916 644702 437994 644802
rect 438118 644702 438218 644802
rect 438342 644702 438442 644802
rect 438566 644702 438666 644802
rect 438790 644702 438890 644802
rect 437894 644478 437916 644578
rect 437916 644478 437994 644578
rect 438118 644478 438218 644578
rect 438342 644478 438442 644578
rect 438566 644478 438666 644578
rect 438790 644478 438890 644578
rect 437894 644254 437916 644354
rect 437916 644254 437994 644354
rect 438118 644254 438218 644354
rect 438342 644254 438442 644354
rect 438566 644254 438666 644354
rect 438790 644254 438890 644354
rect 437894 644030 437916 644130
rect 437916 644030 437994 644130
rect 438118 644030 438218 644130
rect 438342 644030 438442 644130
rect 438566 644030 438666 644130
rect 438790 644030 438890 644130
rect 437894 643806 437916 643906
rect 437916 643806 437994 643906
rect 438118 643806 438218 643906
rect 438342 643806 438442 643906
rect 438566 643806 438666 643906
rect 438790 643806 438890 643906
rect 437894 643582 437916 643682
rect 437916 643582 437994 643682
rect 438118 643582 438218 643682
rect 438342 643582 438442 643682
rect 438566 643582 438666 643682
rect 438790 643582 438890 643682
rect 437894 636678 437916 636778
rect 437916 636678 437994 636778
rect 438118 636678 438218 636778
rect 438342 636678 438442 636778
rect 438566 636678 438666 636778
rect 438790 636678 438890 636778
rect 437894 636454 437916 636554
rect 437916 636454 437994 636554
rect 438118 636454 438218 636554
rect 438342 636454 438442 636554
rect 438566 636454 438666 636554
rect 438790 636454 438890 636554
rect 437894 636230 437916 636330
rect 437916 636230 437994 636330
rect 438118 636230 438218 636330
rect 438342 636230 438442 636330
rect 438566 636230 438666 636330
rect 438790 636230 438890 636330
rect 437894 636006 437916 636106
rect 437916 636006 437994 636106
rect 438118 636006 438218 636106
rect 438342 636006 438442 636106
rect 438566 636006 438666 636106
rect 438790 636006 438890 636106
rect 437894 635782 437916 635882
rect 437916 635782 437994 635882
rect 438118 635782 438218 635882
rect 438342 635782 438442 635882
rect 438566 635782 438666 635882
rect 438790 635782 438890 635882
rect 437894 635558 437916 635658
rect 437916 635558 437994 635658
rect 438118 635558 438218 635658
rect 438342 635558 438442 635658
rect 438566 635558 438666 635658
rect 438790 635558 438890 635658
rect 437894 635334 437916 635434
rect 437916 635334 437994 635434
rect 438118 635334 438218 635434
rect 438342 635334 438442 635434
rect 438566 635334 438666 635434
rect 438790 635334 438890 635434
rect 437894 635110 437916 635210
rect 437916 635110 437994 635210
rect 438118 635110 438218 635210
rect 438342 635110 438442 635210
rect 438566 635110 438666 635210
rect 438790 635110 438890 635210
rect 437894 634886 437916 634986
rect 437916 634886 437994 634986
rect 438118 634886 438218 634986
rect 438342 634886 438442 634986
rect 438566 634886 438666 634986
rect 438790 634886 438890 634986
rect 437894 634662 437916 634762
rect 437916 634662 437994 634762
rect 438118 634662 438218 634762
rect 438342 634662 438442 634762
rect 438566 634662 438666 634762
rect 438790 634662 438890 634762
rect 437894 634438 437916 634538
rect 437916 634438 437994 634538
rect 438118 634438 438218 634538
rect 438342 634438 438442 634538
rect 438566 634438 438666 634538
rect 438790 634438 438890 634538
rect 437894 634214 437916 634314
rect 437916 634214 437994 634314
rect 438118 634214 438218 634314
rect 438342 634214 438442 634314
rect 438566 634214 438666 634314
rect 438790 634214 438890 634314
rect 437894 633990 437916 634090
rect 437916 633990 437994 634090
rect 438118 633990 438218 634090
rect 438342 633990 438442 634090
rect 438566 633990 438666 634090
rect 438790 633990 438890 634090
rect 437894 633766 437916 633866
rect 437916 633766 437994 633866
rect 438118 633766 438218 633866
rect 438342 633766 438442 633866
rect 438566 633766 438666 633866
rect 438790 633766 438890 633866
rect 437894 633542 437916 633642
rect 437916 633542 437994 633642
rect 438118 633542 438218 633642
rect 438342 633542 438442 633642
rect 438566 633542 438666 633642
rect 438790 633542 438890 633642
rect 437894 633318 437916 633418
rect 437916 633318 437994 633418
rect 438118 633318 438218 633418
rect 438342 633318 438442 633418
rect 438566 633318 438666 633418
rect 438790 633318 438890 633418
rect 437894 633094 437916 633194
rect 437916 633094 437994 633194
rect 438118 633094 438218 633194
rect 438342 633094 438442 633194
rect 438566 633094 438666 633194
rect 438790 633094 438890 633194
rect 437894 632870 437916 632970
rect 437916 632870 437994 632970
rect 438118 632870 438218 632970
rect 438342 632870 438442 632970
rect 438566 632870 438666 632970
rect 438790 632870 438890 632970
rect 437894 632646 437916 632746
rect 437916 632646 437994 632746
rect 438118 632646 438218 632746
rect 438342 632646 438442 632746
rect 438566 632646 438666 632746
rect 438790 632646 438890 632746
rect 437894 632422 437916 632522
rect 437916 632422 437994 632522
rect 438118 632422 438218 632522
rect 438342 632422 438442 632522
rect 438566 632422 438666 632522
rect 438790 632422 438890 632522
rect 437894 632198 437916 632298
rect 437916 632198 437994 632298
rect 438118 632198 438218 632298
rect 438342 632198 438442 632298
rect 438566 632198 438666 632298
rect 438790 632198 438890 632298
rect 437894 631974 437916 632074
rect 437916 631974 437994 632074
rect 438118 631974 438218 632074
rect 438342 631974 438442 632074
rect 438566 631974 438666 632074
rect 438790 631974 438890 632074
rect 437894 631750 437916 631850
rect 437916 631750 437994 631850
rect 438118 631750 438218 631850
rect 438342 631750 438442 631850
rect 438566 631750 438666 631850
rect 438790 631750 438890 631850
rect 437894 631526 437916 631626
rect 437916 631526 437994 631626
rect 438118 631526 438218 631626
rect 438342 631526 438442 631626
rect 438566 631526 438666 631626
rect 438790 631526 438890 631626
rect 437894 631302 437916 631402
rect 437916 631302 437994 631402
rect 438118 631302 438218 631402
rect 438342 631302 438442 631402
rect 438566 631302 438666 631402
rect 438790 631302 438890 631402
rect 437894 631078 437916 631178
rect 437916 631078 437994 631178
rect 438118 631078 438218 631178
rect 438342 631078 438442 631178
rect 438566 631078 438666 631178
rect 438790 631078 438890 631178
rect 437894 630854 437916 630954
rect 437916 630854 437994 630954
rect 438118 630854 438218 630954
rect 438342 630854 438442 630954
rect 438566 630854 438666 630954
rect 438790 630854 438890 630954
rect 437894 630630 437916 630730
rect 437916 630630 437994 630730
rect 438118 630630 438218 630730
rect 438342 630630 438442 630730
rect 438566 630630 438666 630730
rect 438790 630630 438890 630730
rect 437894 630406 437916 630506
rect 437916 630406 437994 630506
rect 438118 630406 438218 630506
rect 438342 630406 438442 630506
rect 438566 630406 438666 630506
rect 438790 630406 438890 630506
rect 437894 630182 437916 630282
rect 437916 630182 437994 630282
rect 438118 630182 438218 630282
rect 438342 630182 438442 630282
rect 438566 630182 438666 630282
rect 438790 630182 438890 630282
rect 440716 652724 451932 652740
rect 440716 651958 440732 652724
rect 440732 651958 451916 652724
rect 451916 651958 451932 652724
rect 440716 651942 451932 651958
rect 456604 649267 457142 649664
rect 457422 649267 457960 649664
rect 458240 649267 458778 649664
rect 459058 649267 459596 649664
rect 461512 649205 462050 649602
rect 462330 649205 462868 649602
rect 463148 649205 463686 649602
rect 463966 649205 464504 649602
rect 464784 649205 465322 649602
rect 465602 649205 466140 649602
rect 466420 649205 466958 649602
rect 467238 649205 467776 649602
rect 468056 649205 468594 649602
rect 468874 649205 469412 649602
rect 469692 649205 470230 649602
rect 470510 649205 471048 649602
rect 471328 649205 471866 649602
rect 472146 649205 472684 649602
rect 472964 649205 473502 649602
rect 473782 649205 474320 649602
rect 474600 649205 475138 649602
rect 453332 647881 453870 648278
rect 454150 647881 454688 648278
rect 454968 647881 455506 648278
rect 453332 644126 453870 644523
rect 454150 644126 454688 644523
rect 454968 644126 455506 644523
rect 455788 643856 456282 644922
rect 456604 644536 457142 644933
rect 457422 644536 457960 644933
rect 458240 644536 458778 644933
rect 459058 644536 459596 644933
rect 460740 643868 461252 644920
rect 461512 642470 462050 642867
rect 462330 642469 462868 642867
rect 463148 642470 463686 642867
rect 463966 642470 464504 642867
rect 464784 642469 465322 642867
rect 465602 642470 466140 642867
rect 466420 642470 466958 642867
rect 467238 642469 467776 642867
rect 468056 642470 468594 642867
rect 468874 642470 469412 642867
rect 469692 642470 470230 642867
rect 470510 642469 471048 642867
rect 471328 642470 471866 642867
rect 472146 642470 472684 642867
rect 472964 642470 473502 642867
rect 473782 642470 474320 642867
rect 474600 642470 475138 642867
rect 444360 637070 450824 637076
rect 444360 636738 444366 637070
rect 444366 636738 450818 637070
rect 450818 636738 450824 637070
rect 444360 636732 450824 636738
rect 445084 636506 450460 636540
rect 445000 636202 445034 636386
rect 445084 636048 450460 636082
rect 445520 634380 445704 634414
rect 446092 634380 446276 634414
rect 446664 634380 446848 634414
rect 447236 634380 447420 634414
rect 447808 634380 447992 634414
rect 448380 634380 448564 634414
rect 448952 634380 449136 634414
rect 449524 634380 449708 634414
rect 441342 633356 441394 633408
rect 442258 633356 442310 633408
rect 440590 633258 440774 633292
rect 441048 633258 441232 633292
rect 441506 633258 441690 633292
rect 441964 633258 442148 633292
rect 442422 633258 442606 633292
rect 442880 633258 443064 633292
rect 440436 632832 440470 633208
rect 440894 632832 440928 633208
rect 441352 632832 441386 633208
rect 441810 632832 441844 633208
rect 442268 632832 442302 633208
rect 442726 632832 442760 633208
rect 443184 632832 443218 633208
rect 444814 632732 444914 634330
rect 445366 632554 445400 634330
rect 445824 632554 445858 634330
rect 445938 632554 445972 634330
rect 446396 632554 446430 634330
rect 446510 632554 446544 634330
rect 446968 632554 447002 634330
rect 447082 632554 447116 634330
rect 447540 632554 447574 634330
rect 447654 632554 447688 634330
rect 448112 632554 448146 634330
rect 448226 632554 448260 634330
rect 448684 632554 448718 634330
rect 448798 632554 448832 634330
rect 449256 632554 449290 634330
rect 449370 632554 449404 634330
rect 449828 632554 449862 634330
rect 450314 632732 450414 634330
rect 443794 631977 443978 632011
rect 444366 631977 444550 632011
rect 444938 631977 445122 632011
rect 445510 631977 445694 632011
rect 446082 631977 446266 632011
rect 446654 631977 446838 632011
rect 447226 631977 447410 632011
rect 447798 631977 447982 632011
rect 448370 631977 448554 632011
rect 448942 631977 449126 632011
rect 449514 631977 449698 632011
rect 450086 631977 450270 632011
rect 450658 631977 450842 632011
rect 451230 631977 451414 632011
rect 442998 629488 443098 631830
rect 443640 629362 443674 631918
rect 444098 629362 444132 631918
rect 444212 629362 444246 631918
rect 444670 629362 444704 631918
rect 444784 629362 444818 631918
rect 445242 629362 445276 631918
rect 445356 629362 445390 631918
rect 445814 629362 445848 631918
rect 445928 629362 445962 631918
rect 446386 629362 446420 631918
rect 446500 629362 446534 631918
rect 446958 629362 446992 631918
rect 447072 629362 447106 631918
rect 447530 629362 447564 631918
rect 447644 629362 447678 631918
rect 448102 629362 448136 631918
rect 448216 629362 448250 631918
rect 448674 629362 448708 631918
rect 448788 629362 448822 631918
rect 449246 629362 449280 631918
rect 449360 629362 449394 631918
rect 449818 629362 449852 631918
rect 449932 629362 449966 631918
rect 450390 629362 450424 631918
rect 450504 629362 450538 631918
rect 450962 629362 450996 631918
rect 451076 629362 451110 631918
rect 451534 629362 451568 631918
rect 452126 629488 452226 631830
rect 446580 628884 448922 628984
rect 453448 629400 453482 637116
rect 453906 629400 453940 637116
rect 454364 629400 454398 637116
rect 454822 629400 454856 637116
rect 455280 629400 455314 637116
rect 455738 629400 455772 637116
rect 456196 629400 456230 637116
rect 456654 629400 456688 637116
rect 457112 629400 457146 637116
rect 457570 629400 457604 637116
rect 458028 629400 458062 637116
rect 458486 629400 458520 637116
rect 453602 629307 453786 629341
rect 454060 629307 454244 629341
rect 454518 629307 454702 629341
rect 454976 629307 455160 629341
rect 455434 629307 455618 629341
rect 455892 629307 456076 629341
rect 456350 629307 456534 629341
rect 456808 629307 456992 629341
rect 457266 629307 457450 629341
rect 457724 629307 457908 629341
rect 458182 629307 458366 629341
rect 452848 628790 453248 628890
rect 459406 629400 459440 637116
rect 459864 629400 459898 637116
rect 460322 629400 460356 637116
rect 460780 629400 460814 637116
rect 461238 629400 461272 637116
rect 461696 629400 461730 637116
rect 462154 629400 462188 637116
rect 462612 629400 462646 637116
rect 463070 629400 463104 637116
rect 463528 629400 463562 637116
rect 463986 629400 464020 637116
rect 459560 629307 459744 629341
rect 460018 629307 460202 629341
rect 460476 629307 460660 629341
rect 460934 629307 461118 629341
rect 461392 629307 461576 629341
rect 461850 629307 462034 629341
rect 462308 629307 462492 629341
rect 462766 629307 462950 629341
rect 463224 629307 463408 629341
rect 463682 629307 463866 629341
rect 458758 628790 459158 628890
rect 464906 629400 464940 637116
rect 465364 629400 465398 637116
rect 465822 629400 465856 637116
rect 466280 629400 466314 637116
rect 466738 629400 466772 637116
rect 467196 629400 467230 637116
rect 467654 629400 467688 637116
rect 468112 629400 468146 637116
rect 468570 629400 468604 637116
rect 469028 629400 469062 637116
rect 469486 629400 469520 637116
rect 469944 629400 469978 637116
rect 465060 629307 465244 629341
rect 465518 629307 465702 629341
rect 465976 629307 466160 629341
rect 466434 629307 466618 629341
rect 466892 629307 467076 629341
rect 467350 629307 467534 629341
rect 467808 629307 467992 629341
rect 468266 629307 468450 629341
rect 468724 629307 468908 629341
rect 469182 629307 469366 629341
rect 469640 629307 469824 629341
rect 464258 628790 464658 628890
rect 470214 628788 470614 628888
rect 438920 627630 439020 627656
rect 439144 627630 439244 627656
rect 439368 627630 439468 627656
rect 439592 627630 439692 627656
rect 439816 627630 439916 627656
rect 440040 627630 440140 627656
rect 440264 627630 440364 627656
rect 440488 627630 440588 627656
rect 440712 627630 440812 627656
rect 440936 627630 441036 627656
rect 441160 627630 441260 627656
rect 441384 627630 441484 627656
rect 441608 627630 441708 627656
rect 441832 627630 441932 627656
rect 442056 627630 442156 627656
rect 442280 627630 442380 627656
rect 442504 627630 442604 627656
rect 442728 627630 442828 627656
rect 442952 627630 443052 627656
rect 443176 627630 443276 627656
rect 443400 627630 443500 627656
rect 443624 627630 443724 627656
rect 443848 627630 443948 627656
rect 444072 627630 444172 627656
rect 444296 627630 444396 627656
rect 444520 627630 444620 627656
rect 444744 627630 444844 627656
rect 444968 627630 445068 627656
rect 445192 627630 445292 627656
rect 445416 627630 445516 627656
rect 449390 627630 449490 627656
rect 449614 627630 449714 627656
rect 449838 627630 449938 627656
rect 450062 627630 450162 627656
rect 450286 627630 450386 627656
rect 450510 627630 450610 627656
rect 450734 627630 450834 627656
rect 450958 627630 451058 627656
rect 451182 627630 451282 627656
rect 451406 627630 451506 627656
rect 451630 627630 451730 627656
rect 451854 627630 451954 627656
rect 452078 627630 452178 627656
rect 452302 627630 452402 627656
rect 452526 627630 452626 627656
rect 452750 627630 452850 627656
rect 452974 627630 453074 627656
rect 453198 627630 453298 627656
rect 453422 627630 453522 627656
rect 453646 627630 453746 627656
rect 453870 627630 453970 627656
rect 454094 627630 454194 627656
rect 454318 627630 454418 627656
rect 454542 627630 454642 627656
rect 454766 627630 454866 627656
rect 454990 627630 455090 627656
rect 455214 627630 455314 627656
rect 455438 627630 455538 627656
rect 455662 627630 455762 627656
rect 455886 627630 455986 627656
rect 475660 627630 475760 627676
rect 475884 627630 475984 627676
rect 476108 627630 476208 627676
rect 476332 627630 476432 627676
rect 476556 627630 476656 627676
rect 476780 627630 476880 627676
rect 477004 627630 477104 627676
rect 477228 627630 477328 627676
rect 477452 627630 477552 627676
rect 477676 627630 477776 627676
rect 477900 627630 478000 627676
rect 478124 627630 478224 627676
rect 478348 627630 478448 627676
rect 478572 627630 478672 627676
rect 478796 627630 478896 627676
rect 479020 627630 479120 627676
rect 479244 627630 479344 627676
rect 479468 627630 479568 627676
rect 479692 627630 479792 627676
rect 479916 627630 480016 627676
rect 480140 627630 480240 627676
rect 480364 627630 480464 627676
rect 480588 627630 480688 627676
rect 480812 627630 480912 627676
rect 481036 627630 481136 627676
rect 438920 627556 439020 627630
rect 439144 627556 439244 627630
rect 439368 627556 439468 627630
rect 439592 627556 439692 627630
rect 439816 627556 439916 627630
rect 440040 627556 440140 627630
rect 440264 627556 440364 627630
rect 440488 627556 440588 627630
rect 440712 627556 440812 627630
rect 440936 627556 441036 627630
rect 441160 627556 441260 627630
rect 441384 627556 441484 627630
rect 441608 627556 441708 627630
rect 441832 627556 441932 627630
rect 442056 627556 442156 627630
rect 442280 627556 442380 627630
rect 442504 627556 442604 627630
rect 442728 627556 442828 627630
rect 442952 627556 443052 627630
rect 443176 627556 443276 627630
rect 443400 627556 443500 627630
rect 443624 627556 443724 627630
rect 443848 627556 443948 627630
rect 444072 627556 444172 627630
rect 444296 627556 444396 627630
rect 444520 627556 444620 627630
rect 444744 627556 444844 627630
rect 444968 627556 445068 627630
rect 445192 627556 445292 627630
rect 445416 627556 445516 627630
rect 449390 627556 449490 627630
rect 449614 627556 449714 627630
rect 449838 627556 449938 627630
rect 450062 627556 450162 627630
rect 450286 627556 450386 627630
rect 450510 627556 450610 627630
rect 450734 627556 450834 627630
rect 450958 627556 451058 627630
rect 451182 627556 451282 627630
rect 451406 627556 451506 627630
rect 451630 627556 451730 627630
rect 451854 627556 451954 627630
rect 452078 627556 452178 627630
rect 452302 627556 452402 627630
rect 452526 627556 452626 627630
rect 452750 627556 452850 627630
rect 452974 627556 453074 627630
rect 453198 627556 453298 627630
rect 453422 627556 453522 627630
rect 453646 627556 453746 627630
rect 453870 627556 453970 627630
rect 454094 627556 454194 627630
rect 454318 627556 454418 627630
rect 454542 627556 454642 627630
rect 454766 627556 454866 627630
rect 454990 627556 455090 627630
rect 455214 627556 455314 627630
rect 455438 627556 455538 627630
rect 455662 627556 455762 627630
rect 455886 627556 455986 627630
rect 475660 627576 475760 627630
rect 475884 627576 475984 627630
rect 476108 627576 476208 627630
rect 476332 627576 476432 627630
rect 476556 627576 476656 627630
rect 476780 627576 476880 627630
rect 477004 627576 477104 627630
rect 477228 627576 477328 627630
rect 477452 627576 477552 627630
rect 477676 627576 477776 627630
rect 477900 627576 478000 627630
rect 478124 627576 478224 627630
rect 478348 627576 478448 627630
rect 478572 627576 478672 627630
rect 478796 627576 478896 627630
rect 479020 627576 479120 627630
rect 479244 627576 479344 627630
rect 479468 627576 479568 627630
rect 479692 627576 479792 627630
rect 479916 627576 480016 627630
rect 480140 627576 480240 627630
rect 480364 627576 480464 627630
rect 480588 627576 480688 627630
rect 480812 627576 480912 627630
rect 481036 627576 481132 627630
rect 481132 627576 481136 627630
rect 481260 627576 481360 627676
rect 481484 627576 481584 627676
rect 481708 627576 481808 627676
rect 481932 627576 482032 627676
rect 482174 650078 482274 650178
rect 482398 650078 482498 650178
rect 482622 650078 482722 650178
rect 482846 650078 482946 650178
rect 483070 650078 483156 650178
rect 483156 650078 483170 650178
rect 482174 649854 482274 649954
rect 482398 649854 482498 649954
rect 482622 649854 482722 649954
rect 482846 649854 482946 649954
rect 483070 649854 483156 649954
rect 483156 649854 483170 649954
rect 482174 649630 482274 649730
rect 482398 649630 482498 649730
rect 482622 649630 482722 649730
rect 482846 649630 482946 649730
rect 483070 649630 483156 649730
rect 483156 649630 483170 649730
rect 482174 649406 482274 649506
rect 482398 649406 482498 649506
rect 482622 649406 482722 649506
rect 482846 649406 482946 649506
rect 483070 649406 483156 649506
rect 483156 649406 483170 649506
rect 482174 649182 482274 649282
rect 482398 649182 482498 649282
rect 482622 649182 482722 649282
rect 482846 649182 482946 649282
rect 483070 649182 483156 649282
rect 483156 649182 483170 649282
rect 482174 648958 482274 649058
rect 482398 648958 482498 649058
rect 482622 648958 482722 649058
rect 482846 648958 482946 649058
rect 483070 648958 483156 649058
rect 483156 648958 483170 649058
rect 482174 648734 482274 648834
rect 482398 648734 482498 648834
rect 482622 648734 482722 648834
rect 482846 648734 482946 648834
rect 483070 648734 483156 648834
rect 483156 648734 483170 648834
rect 482174 648510 482274 648610
rect 482398 648510 482498 648610
rect 482622 648510 482722 648610
rect 482846 648510 482946 648610
rect 483070 648510 483156 648610
rect 483156 648510 483170 648610
rect 482174 648286 482274 648386
rect 482398 648286 482498 648386
rect 482622 648286 482722 648386
rect 482846 648286 482946 648386
rect 483070 648286 483156 648386
rect 483156 648286 483170 648386
rect 482174 648062 482274 648162
rect 482398 648062 482498 648162
rect 482622 648062 482722 648162
rect 482846 648062 482946 648162
rect 483070 648062 483156 648162
rect 483156 648062 483170 648162
rect 482174 647838 482274 647938
rect 482398 647838 482498 647938
rect 482622 647838 482722 647938
rect 482846 647838 482946 647938
rect 483070 647838 483156 647938
rect 483156 647838 483170 647938
rect 482174 647614 482274 647714
rect 482398 647614 482498 647714
rect 482622 647614 482722 647714
rect 482846 647614 482946 647714
rect 483070 647614 483156 647714
rect 483156 647614 483170 647714
rect 482174 647390 482274 647490
rect 482398 647390 482498 647490
rect 482622 647390 482722 647490
rect 482846 647390 482946 647490
rect 483070 647390 483156 647490
rect 483156 647390 483170 647490
rect 482174 647166 482274 647266
rect 482398 647166 482498 647266
rect 482622 647166 482722 647266
rect 482846 647166 482946 647266
rect 483070 647166 483156 647266
rect 483156 647166 483170 647266
rect 482174 646942 482274 647042
rect 482398 646942 482498 647042
rect 482622 646942 482722 647042
rect 482846 646942 482946 647042
rect 483070 646942 483156 647042
rect 483156 646942 483170 647042
rect 482174 646718 482274 646818
rect 482398 646718 482498 646818
rect 482622 646718 482722 646818
rect 482846 646718 482946 646818
rect 483070 646718 483156 646818
rect 483156 646718 483170 646818
rect 482174 646494 482274 646594
rect 482398 646494 482498 646594
rect 482622 646494 482722 646594
rect 482846 646494 482946 646594
rect 483070 646494 483156 646594
rect 483156 646494 483170 646594
rect 482174 646270 482274 646370
rect 482398 646270 482498 646370
rect 482622 646270 482722 646370
rect 482846 646270 482946 646370
rect 483070 646270 483156 646370
rect 483156 646270 483170 646370
rect 482174 646046 482274 646146
rect 482398 646046 482498 646146
rect 482622 646046 482722 646146
rect 482846 646046 482946 646146
rect 483070 646046 483156 646146
rect 483156 646046 483170 646146
rect 482174 645822 482274 645922
rect 482398 645822 482498 645922
rect 482622 645822 482722 645922
rect 482846 645822 482946 645922
rect 483070 645822 483156 645922
rect 483156 645822 483170 645922
rect 482174 645598 482274 645698
rect 482398 645598 482498 645698
rect 482622 645598 482722 645698
rect 482846 645598 482946 645698
rect 483070 645598 483156 645698
rect 483156 645598 483170 645698
rect 482174 645374 482274 645474
rect 482398 645374 482498 645474
rect 482622 645374 482722 645474
rect 482846 645374 482946 645474
rect 483070 645374 483156 645474
rect 483156 645374 483170 645474
rect 482174 645150 482274 645250
rect 482398 645150 482498 645250
rect 482622 645150 482722 645250
rect 482846 645150 482946 645250
rect 483070 645150 483156 645250
rect 483156 645150 483170 645250
rect 482174 644926 482274 645026
rect 482398 644926 482498 645026
rect 482622 644926 482722 645026
rect 482846 644926 482946 645026
rect 483070 644926 483156 645026
rect 483156 644926 483170 645026
rect 482174 644702 482274 644802
rect 482398 644702 482498 644802
rect 482622 644702 482722 644802
rect 482846 644702 482946 644802
rect 483070 644702 483156 644802
rect 483156 644702 483170 644802
rect 482174 644478 482274 644578
rect 482398 644478 482498 644578
rect 482622 644478 482722 644578
rect 482846 644478 482946 644578
rect 483070 644478 483156 644578
rect 483156 644478 483170 644578
rect 482174 644254 482274 644354
rect 482398 644254 482498 644354
rect 482622 644254 482722 644354
rect 482846 644254 482946 644354
rect 483070 644254 483156 644354
rect 483156 644254 483170 644354
rect 482174 644030 482274 644130
rect 482398 644030 482498 644130
rect 482622 644030 482722 644130
rect 482846 644030 482946 644130
rect 483070 644030 483156 644130
rect 483156 644030 483170 644130
rect 482174 643806 482274 643906
rect 482398 643806 482498 643906
rect 482622 643806 482722 643906
rect 482846 643806 482946 643906
rect 483070 643806 483156 643906
rect 483156 643806 483170 643906
rect 482174 643582 482274 643682
rect 482398 643582 482498 643682
rect 482622 643582 482722 643682
rect 482846 643582 482946 643682
rect 483070 643582 483156 643682
rect 483156 643582 483170 643682
rect 482174 636678 482274 636778
rect 482398 636678 482498 636778
rect 482622 636678 482722 636778
rect 482846 636678 482946 636778
rect 483070 636678 483156 636778
rect 483156 636678 483170 636778
rect 482174 636454 482274 636554
rect 482398 636454 482498 636554
rect 482622 636454 482722 636554
rect 482846 636454 482946 636554
rect 483070 636454 483156 636554
rect 483156 636454 483170 636554
rect 482174 636230 482274 636330
rect 482398 636230 482498 636330
rect 482622 636230 482722 636330
rect 482846 636230 482946 636330
rect 483070 636230 483156 636330
rect 483156 636230 483170 636330
rect 482174 636006 482274 636106
rect 482398 636006 482498 636106
rect 482622 636006 482722 636106
rect 482846 636006 482946 636106
rect 483070 636006 483156 636106
rect 483156 636006 483170 636106
rect 482174 635782 482274 635882
rect 482398 635782 482498 635882
rect 482622 635782 482722 635882
rect 482846 635782 482946 635882
rect 483070 635782 483156 635882
rect 483156 635782 483170 635882
rect 482174 635558 482274 635658
rect 482398 635558 482498 635658
rect 482622 635558 482722 635658
rect 482846 635558 482946 635658
rect 483070 635558 483156 635658
rect 483156 635558 483170 635658
rect 482174 635334 482274 635434
rect 482398 635334 482498 635434
rect 482622 635334 482722 635434
rect 482846 635334 482946 635434
rect 483070 635334 483156 635434
rect 483156 635334 483170 635434
rect 482174 635110 482274 635210
rect 482398 635110 482498 635210
rect 482622 635110 482722 635210
rect 482846 635110 482946 635210
rect 483070 635110 483156 635210
rect 483156 635110 483170 635210
rect 482174 634886 482274 634986
rect 482398 634886 482498 634986
rect 482622 634886 482722 634986
rect 482846 634886 482946 634986
rect 483070 634886 483156 634986
rect 483156 634886 483170 634986
rect 482174 634662 482274 634762
rect 482398 634662 482498 634762
rect 482622 634662 482722 634762
rect 482846 634662 482946 634762
rect 483070 634662 483156 634762
rect 483156 634662 483170 634762
rect 482174 634438 482274 634538
rect 482398 634438 482498 634538
rect 482622 634438 482722 634538
rect 482846 634438 482946 634538
rect 483070 634438 483156 634538
rect 483156 634438 483170 634538
rect 482174 634214 482274 634314
rect 482398 634214 482498 634314
rect 482622 634214 482722 634314
rect 482846 634214 482946 634314
rect 483070 634214 483156 634314
rect 483156 634214 483170 634314
rect 482174 633990 482274 634090
rect 482398 633990 482498 634090
rect 482622 633990 482722 634090
rect 482846 633990 482946 634090
rect 483070 633990 483156 634090
rect 483156 633990 483170 634090
rect 482174 633766 482274 633866
rect 482398 633766 482498 633866
rect 482622 633766 482722 633866
rect 482846 633766 482946 633866
rect 483070 633766 483156 633866
rect 483156 633766 483170 633866
rect 482174 633542 482274 633642
rect 482398 633542 482498 633642
rect 482622 633542 482722 633642
rect 482846 633542 482946 633642
rect 483070 633542 483156 633642
rect 483156 633542 483170 633642
rect 482174 633318 482274 633418
rect 482398 633318 482498 633418
rect 482622 633318 482722 633418
rect 482846 633318 482946 633418
rect 483070 633318 483156 633418
rect 483156 633318 483170 633418
rect 482174 633094 482274 633194
rect 482398 633094 482498 633194
rect 482622 633094 482722 633194
rect 482846 633094 482946 633194
rect 483070 633094 483156 633194
rect 483156 633094 483170 633194
rect 482174 632870 482274 632970
rect 482398 632870 482498 632970
rect 482622 632870 482722 632970
rect 482846 632870 482946 632970
rect 483070 632870 483156 632970
rect 483156 632870 483170 632970
rect 482174 632646 482274 632746
rect 482398 632646 482498 632746
rect 482622 632646 482722 632746
rect 482846 632646 482946 632746
rect 483070 632646 483156 632746
rect 483156 632646 483170 632746
rect 482174 632422 482274 632522
rect 482398 632422 482498 632522
rect 482622 632422 482722 632522
rect 482846 632422 482946 632522
rect 483070 632422 483156 632522
rect 483156 632422 483170 632522
rect 482174 632198 482274 632298
rect 482398 632198 482498 632298
rect 482622 632198 482722 632298
rect 482846 632198 482946 632298
rect 483070 632198 483156 632298
rect 483156 632198 483170 632298
rect 482174 631974 482274 632074
rect 482398 631974 482498 632074
rect 482622 631974 482722 632074
rect 482846 631974 482946 632074
rect 483070 631974 483156 632074
rect 483156 631974 483170 632074
rect 482174 631750 482274 631850
rect 482398 631750 482498 631850
rect 482622 631750 482722 631850
rect 482846 631750 482946 631850
rect 483070 631750 483156 631850
rect 483156 631750 483170 631850
rect 482174 631526 482274 631626
rect 482398 631526 482498 631626
rect 482622 631526 482722 631626
rect 482846 631526 482946 631626
rect 483070 631526 483156 631626
rect 483156 631526 483170 631626
rect 482174 631302 482274 631402
rect 482398 631302 482498 631402
rect 482622 631302 482722 631402
rect 482846 631302 482946 631402
rect 483070 631302 483156 631402
rect 483156 631302 483170 631402
rect 482174 631078 482274 631178
rect 482398 631078 482498 631178
rect 482622 631078 482722 631178
rect 482846 631078 482946 631178
rect 483070 631078 483156 631178
rect 483156 631078 483170 631178
rect 482174 630854 482274 630954
rect 482398 630854 482498 630954
rect 482622 630854 482722 630954
rect 482846 630854 482946 630954
rect 483070 630854 483156 630954
rect 483156 630854 483170 630954
rect 482174 630630 482274 630730
rect 482398 630630 482498 630730
rect 482622 630630 482722 630730
rect 482846 630630 482946 630730
rect 483070 630630 483156 630730
rect 483156 630630 483170 630730
rect 482174 630406 482274 630506
rect 482398 630406 482498 630506
rect 482622 630406 482722 630506
rect 482846 630406 482946 630506
rect 483070 630406 483156 630506
rect 483156 630406 483170 630506
rect 482174 630182 482274 630282
rect 482398 630182 482498 630282
rect 482622 630182 482722 630282
rect 482846 630182 482946 630282
rect 483070 630182 483156 630282
rect 483156 630182 483170 630282
rect 482156 627576 482256 627676
rect 438920 627332 439020 627432
rect 439144 627332 439244 627432
rect 439368 627332 439468 627432
rect 439592 627332 439692 627432
rect 439816 627332 439916 627432
rect 440040 627332 440140 627432
rect 440264 627332 440364 627432
rect 440488 627332 440588 627432
rect 440712 627332 440812 627432
rect 440936 627332 441036 627432
rect 441160 627332 441260 627432
rect 441384 627332 441484 627432
rect 441608 627332 441708 627432
rect 441832 627332 441932 627432
rect 442056 627332 442156 627432
rect 442280 627332 442380 627432
rect 442504 627332 442604 627432
rect 442728 627332 442828 627432
rect 442952 627332 443052 627432
rect 443176 627332 443276 627432
rect 443400 627332 443500 627432
rect 443624 627332 443724 627432
rect 443848 627332 443948 627432
rect 444072 627332 444172 627432
rect 444296 627332 444396 627432
rect 444520 627332 444620 627432
rect 444744 627332 444844 627432
rect 444968 627332 445068 627432
rect 445192 627332 445292 627432
rect 445416 627332 445516 627432
rect 449390 627332 449490 627432
rect 449614 627332 449714 627432
rect 449838 627332 449938 627432
rect 450062 627332 450162 627432
rect 450286 627332 450386 627432
rect 450510 627332 450610 627432
rect 450734 627332 450834 627432
rect 450958 627332 451058 627432
rect 451182 627332 451282 627432
rect 451406 627332 451506 627432
rect 451630 627332 451730 627432
rect 451854 627332 451954 627432
rect 452078 627332 452178 627432
rect 452302 627332 452402 627432
rect 452526 627332 452626 627432
rect 452750 627332 452850 627432
rect 452974 627332 453074 627432
rect 453198 627332 453298 627432
rect 453422 627332 453522 627432
rect 453646 627332 453746 627432
rect 453870 627332 453970 627432
rect 454094 627332 454194 627432
rect 454318 627332 454418 627432
rect 454542 627332 454642 627432
rect 454766 627332 454866 627432
rect 454990 627332 455090 627432
rect 455214 627332 455314 627432
rect 455438 627332 455538 627432
rect 455662 627332 455762 627432
rect 455886 627332 455986 627432
rect 475660 627352 475760 627452
rect 475884 627352 475984 627452
rect 476108 627352 476208 627452
rect 476332 627352 476432 627452
rect 476556 627352 476656 627452
rect 476780 627352 476880 627452
rect 477004 627352 477104 627452
rect 477228 627352 477328 627452
rect 477452 627352 477552 627452
rect 477676 627352 477776 627452
rect 477900 627352 478000 627452
rect 478124 627352 478224 627452
rect 478348 627352 478448 627452
rect 478572 627352 478672 627452
rect 478796 627352 478896 627452
rect 479020 627352 479120 627452
rect 479244 627352 479344 627452
rect 479468 627352 479568 627452
rect 479692 627352 479792 627452
rect 479916 627352 480016 627452
rect 480140 627352 480240 627452
rect 480364 627352 480464 627452
rect 480588 627352 480688 627452
rect 480812 627352 480912 627452
rect 481036 627352 481132 627452
rect 481132 627352 481136 627452
rect 481260 627352 481360 627452
rect 481484 627352 481584 627452
rect 481708 627352 481808 627452
rect 481932 627352 482032 627452
rect 482156 627352 482256 627452
rect 438920 627108 439020 627208
rect 439144 627108 439244 627208
rect 439368 627108 439468 627208
rect 439592 627108 439692 627208
rect 439816 627108 439916 627208
rect 440040 627108 440140 627208
rect 440264 627108 440364 627208
rect 440488 627108 440588 627208
rect 440712 627108 440812 627208
rect 440936 627108 441036 627208
rect 441160 627108 441260 627208
rect 441384 627108 441484 627208
rect 441608 627108 441708 627208
rect 441832 627108 441932 627208
rect 442056 627108 442156 627208
rect 442280 627108 442380 627208
rect 442504 627108 442604 627208
rect 442728 627108 442828 627208
rect 442952 627108 443052 627208
rect 443176 627108 443276 627208
rect 443400 627108 443500 627208
rect 443624 627108 443724 627208
rect 443848 627108 443948 627208
rect 444072 627108 444172 627208
rect 444296 627108 444396 627208
rect 444520 627108 444620 627208
rect 444744 627108 444844 627208
rect 444968 627108 445068 627208
rect 445192 627108 445292 627208
rect 445416 627108 445516 627208
rect 449390 627108 449490 627208
rect 449614 627108 449714 627208
rect 449838 627108 449938 627208
rect 450062 627108 450162 627208
rect 450286 627108 450386 627208
rect 450510 627108 450610 627208
rect 450734 627108 450834 627208
rect 450958 627108 451058 627208
rect 451182 627108 451282 627208
rect 451406 627108 451506 627208
rect 451630 627108 451730 627208
rect 451854 627108 451954 627208
rect 452078 627108 452178 627208
rect 452302 627108 452402 627208
rect 452526 627108 452626 627208
rect 452750 627108 452850 627208
rect 452974 627108 453074 627208
rect 453198 627108 453298 627208
rect 453422 627108 453522 627208
rect 453646 627108 453746 627208
rect 453870 627108 453970 627208
rect 454094 627108 454194 627208
rect 454318 627108 454418 627208
rect 454542 627108 454642 627208
rect 454766 627108 454866 627208
rect 454990 627108 455090 627208
rect 455214 627108 455314 627208
rect 455438 627108 455538 627208
rect 455662 627108 455762 627208
rect 455886 627108 455986 627208
rect 475660 627128 475760 627228
rect 475884 627128 475984 627228
rect 476108 627128 476208 627228
rect 476332 627128 476432 627228
rect 476556 627128 476656 627228
rect 476780 627128 476880 627228
rect 477004 627128 477104 627228
rect 477228 627128 477328 627228
rect 477452 627128 477552 627228
rect 477676 627128 477776 627228
rect 477900 627128 478000 627228
rect 478124 627128 478224 627228
rect 478348 627128 478448 627228
rect 478572 627128 478672 627228
rect 478796 627128 478896 627228
rect 479020 627128 479120 627228
rect 479244 627128 479344 627228
rect 479468 627128 479568 627228
rect 479692 627128 479792 627228
rect 479916 627128 480016 627228
rect 480140 627128 480240 627228
rect 480364 627128 480464 627228
rect 480588 627128 480688 627228
rect 480812 627128 480912 627228
rect 481036 627128 481132 627228
rect 481132 627128 481136 627228
rect 481260 627128 481360 627228
rect 481484 627128 481584 627228
rect 481708 627128 481808 627228
rect 481932 627128 482032 627228
rect 482156 627128 482256 627228
rect 438920 626884 439020 626984
rect 439144 626884 439244 626984
rect 439368 626884 439468 626984
rect 439592 626884 439692 626984
rect 439816 626884 439916 626984
rect 440040 626884 440140 626984
rect 440264 626884 440364 626984
rect 440488 626884 440588 626984
rect 440712 626884 440812 626984
rect 440936 626884 441036 626984
rect 441160 626884 441260 626984
rect 441384 626884 441484 626984
rect 441608 626884 441708 626984
rect 441832 626884 441932 626984
rect 442056 626884 442156 626984
rect 442280 626884 442380 626984
rect 442504 626884 442604 626984
rect 442728 626884 442828 626984
rect 442952 626884 443052 626984
rect 443176 626884 443276 626984
rect 443400 626884 443500 626984
rect 443624 626884 443724 626984
rect 443848 626884 443948 626984
rect 444072 626884 444172 626984
rect 444296 626884 444396 626984
rect 444520 626884 444620 626984
rect 444744 626884 444844 626984
rect 444968 626884 445068 626984
rect 445192 626884 445292 626984
rect 445416 626884 445516 626984
rect 449390 626884 449490 626984
rect 449614 626884 449714 626984
rect 449838 626884 449938 626984
rect 450062 626884 450162 626984
rect 450286 626884 450386 626984
rect 450510 626884 450610 626984
rect 450734 626884 450834 626984
rect 450958 626884 451058 626984
rect 451182 626884 451282 626984
rect 451406 626884 451506 626984
rect 451630 626884 451730 626984
rect 451854 626884 451954 626984
rect 452078 626884 452178 626984
rect 452302 626884 452402 626984
rect 452526 626884 452626 626984
rect 452750 626884 452850 626984
rect 452974 626884 453074 626984
rect 453198 626884 453298 626984
rect 453422 626884 453522 626984
rect 453646 626884 453746 626984
rect 453870 626884 453970 626984
rect 454094 626884 454194 626984
rect 454318 626884 454418 626984
rect 454542 626884 454642 626984
rect 454766 626884 454866 626984
rect 454990 626884 455090 626984
rect 455214 626884 455314 626984
rect 455438 626884 455538 626984
rect 455662 626884 455762 626984
rect 455886 626884 455986 626984
rect 475660 626904 475760 627004
rect 475884 626904 475984 627004
rect 476108 626904 476208 627004
rect 476332 626904 476432 627004
rect 476556 626904 476656 627004
rect 476780 626904 476880 627004
rect 477004 626904 477104 627004
rect 477228 626904 477328 627004
rect 477452 626904 477552 627004
rect 477676 626904 477776 627004
rect 477900 626904 478000 627004
rect 478124 626904 478224 627004
rect 478348 626904 478448 627004
rect 478572 626904 478672 627004
rect 478796 626904 478896 627004
rect 479020 626904 479120 627004
rect 479244 626904 479344 627004
rect 479468 626904 479568 627004
rect 479692 626904 479792 627004
rect 479916 626904 480016 627004
rect 480140 626904 480240 627004
rect 480364 626904 480464 627004
rect 480588 626904 480688 627004
rect 480812 626904 480912 627004
rect 481036 626904 481132 627004
rect 481132 626904 481136 627004
rect 481260 626904 481360 627004
rect 481484 626904 481584 627004
rect 481708 626904 481808 627004
rect 481932 626904 482032 627004
rect 482156 626904 482256 627004
rect 438920 626660 439020 626760
rect 439144 626660 439244 626760
rect 439368 626660 439468 626760
rect 439592 626660 439692 626760
rect 439816 626660 439916 626760
rect 440040 626660 440140 626760
rect 440264 626660 440364 626760
rect 440488 626660 440588 626760
rect 440712 626660 440812 626760
rect 440936 626660 441036 626760
rect 441160 626660 441260 626760
rect 441384 626660 441484 626760
rect 441608 626660 441708 626760
rect 441832 626660 441932 626760
rect 442056 626660 442156 626760
rect 442280 626660 442380 626760
rect 442504 626660 442604 626760
rect 442728 626660 442828 626760
rect 442952 626660 443052 626760
rect 443176 626660 443276 626760
rect 443400 626660 443500 626760
rect 443624 626660 443724 626760
rect 443848 626660 443948 626760
rect 444072 626660 444172 626760
rect 444296 626660 444396 626760
rect 444520 626660 444620 626760
rect 444744 626660 444844 626760
rect 444968 626660 445068 626760
rect 445192 626660 445292 626760
rect 445416 626660 445516 626760
rect 449390 626660 449490 626760
rect 449614 626660 449714 626760
rect 449838 626660 449938 626760
rect 450062 626660 450162 626760
rect 450286 626660 450386 626760
rect 450510 626660 450610 626760
rect 450734 626660 450834 626760
rect 450958 626660 451058 626760
rect 451182 626660 451282 626760
rect 451406 626660 451506 626760
rect 451630 626660 451730 626760
rect 451854 626660 451954 626760
rect 452078 626660 452178 626760
rect 452302 626660 452402 626760
rect 452526 626660 452626 626760
rect 452750 626660 452850 626760
rect 452974 626660 453074 626760
rect 453198 626660 453298 626760
rect 453422 626660 453522 626760
rect 453646 626660 453746 626760
rect 453870 626660 453970 626760
rect 454094 626660 454194 626760
rect 454318 626660 454418 626760
rect 454542 626660 454642 626760
rect 454766 626660 454866 626760
rect 454990 626660 455090 626760
rect 455214 626660 455314 626760
rect 455438 626660 455538 626760
rect 455662 626660 455762 626760
rect 455886 626660 455986 626760
rect 475660 626680 475760 626780
rect 475884 626680 475984 626780
rect 476108 626680 476208 626780
rect 476332 626680 476432 626780
rect 476556 626680 476656 626780
rect 476780 626680 476880 626780
rect 477004 626680 477104 626780
rect 477228 626680 477328 626780
rect 477452 626680 477552 626780
rect 477676 626680 477776 626780
rect 477900 626680 478000 626780
rect 478124 626680 478224 626780
rect 478348 626680 478448 626780
rect 478572 626680 478672 626780
rect 478796 626680 478896 626780
rect 479020 626680 479120 626780
rect 479244 626680 479344 626780
rect 479468 626680 479568 626780
rect 479692 626680 479792 626780
rect 479916 626680 480016 626780
rect 480140 626680 480240 626780
rect 480364 626680 480464 626780
rect 480588 626680 480688 626780
rect 480812 626680 480912 626780
rect 481036 626680 481132 626780
rect 481132 626680 481136 626780
rect 481260 626680 481360 626780
rect 481484 626680 481584 626780
rect 481708 626680 481808 626780
rect 481932 626680 482032 626780
rect 482156 626680 482256 626780
<< metal1 >>
rect 438880 654876 445540 654906
rect 438880 654776 438920 654876
rect 439020 654776 439144 654876
rect 439244 654776 439368 654876
rect 439468 654776 439592 654876
rect 439692 654776 439816 654876
rect 439916 654776 440040 654876
rect 440140 654776 440264 654876
rect 440364 654776 440488 654876
rect 440588 654776 440712 654876
rect 440812 654776 440936 654876
rect 441036 654776 441160 654876
rect 441260 654776 441384 654876
rect 441484 654776 441608 654876
rect 441708 654776 441832 654876
rect 441932 654776 442056 654876
rect 442156 654776 442280 654876
rect 442380 654776 442504 654876
rect 442604 654776 442728 654876
rect 442828 654776 442952 654876
rect 443052 654776 443176 654876
rect 443276 654776 443400 654876
rect 443500 654776 443624 654876
rect 443724 654776 443848 654876
rect 443948 654776 444072 654876
rect 444172 654776 444296 654876
rect 444396 654776 444520 654876
rect 444620 654776 444744 654876
rect 444844 654776 444968 654876
rect 445068 654776 445192 654876
rect 445292 654776 445416 654876
rect 445516 654776 445540 654876
rect 438880 654652 445540 654776
rect 438880 654552 438920 654652
rect 439020 654552 439144 654652
rect 439244 654552 439368 654652
rect 439468 654552 439592 654652
rect 439692 654552 439816 654652
rect 439916 654552 440040 654652
rect 440140 654552 440264 654652
rect 440364 654552 440488 654652
rect 440588 654552 440712 654652
rect 440812 654552 440936 654652
rect 441036 654552 441160 654652
rect 441260 654552 441384 654652
rect 441484 654552 441608 654652
rect 441708 654552 441832 654652
rect 441932 654552 442056 654652
rect 442156 654552 442280 654652
rect 442380 654552 442504 654652
rect 442604 654552 442728 654652
rect 442828 654552 442952 654652
rect 443052 654552 443176 654652
rect 443276 654552 443400 654652
rect 443500 654552 443624 654652
rect 443724 654552 443848 654652
rect 443948 654552 444072 654652
rect 444172 654552 444296 654652
rect 444396 654552 444520 654652
rect 444620 654552 444744 654652
rect 444844 654552 444968 654652
rect 445068 654552 445192 654652
rect 445292 654552 445416 654652
rect 445516 654552 445540 654652
rect 438880 654428 445540 654552
rect 438880 654328 438920 654428
rect 439020 654328 439144 654428
rect 439244 654328 439368 654428
rect 439468 654328 439592 654428
rect 439692 654328 439816 654428
rect 439916 654328 440040 654428
rect 440140 654328 440264 654428
rect 440364 654328 440488 654428
rect 440588 654328 440712 654428
rect 440812 654328 440936 654428
rect 441036 654328 441160 654428
rect 441260 654328 441384 654428
rect 441484 654328 441608 654428
rect 441708 654328 441832 654428
rect 441932 654328 442056 654428
rect 442156 654328 442280 654428
rect 442380 654328 442504 654428
rect 442604 654328 442728 654428
rect 442828 654328 442952 654428
rect 443052 654328 443176 654428
rect 443276 654328 443400 654428
rect 443500 654328 443624 654428
rect 443724 654328 443848 654428
rect 443948 654328 444072 654428
rect 444172 654328 444296 654428
rect 444396 654328 444520 654428
rect 444620 654328 444744 654428
rect 444844 654328 444968 654428
rect 445068 654328 445192 654428
rect 445292 654328 445416 654428
rect 445516 654328 445540 654428
rect 438880 654204 445540 654328
rect 438880 654104 438920 654204
rect 439020 654104 439144 654204
rect 439244 654104 439368 654204
rect 439468 654104 439592 654204
rect 439692 654104 439816 654204
rect 439916 654104 440040 654204
rect 440140 654104 440264 654204
rect 440364 654104 440488 654204
rect 440588 654104 440712 654204
rect 440812 654104 440936 654204
rect 441036 654104 441160 654204
rect 441260 654104 441384 654204
rect 441484 654104 441608 654204
rect 441708 654104 441832 654204
rect 441932 654104 442056 654204
rect 442156 654104 442280 654204
rect 442380 654104 442504 654204
rect 442604 654104 442728 654204
rect 442828 654104 442952 654204
rect 443052 654104 443176 654204
rect 443276 654104 443400 654204
rect 443500 654104 443624 654204
rect 443724 654104 443848 654204
rect 443948 654104 444072 654204
rect 444172 654104 444296 654204
rect 444396 654104 444520 654204
rect 444620 654104 444744 654204
rect 444844 654104 444968 654204
rect 445068 654104 445192 654204
rect 445292 654104 445416 654204
rect 445516 654104 445540 654204
rect 438880 653980 445540 654104
rect 438880 653880 438920 653980
rect 439020 653880 439144 653980
rect 439244 653880 439368 653980
rect 439468 653880 439592 653980
rect 439692 653880 439816 653980
rect 439916 653880 440040 653980
rect 440140 653880 440264 653980
rect 440364 653880 440488 653980
rect 440588 653880 440712 653980
rect 440812 653880 440936 653980
rect 441036 653880 441160 653980
rect 441260 653880 441384 653980
rect 441484 653880 441608 653980
rect 441708 653880 441832 653980
rect 441932 653880 442056 653980
rect 442156 653880 442280 653980
rect 442380 653880 442504 653980
rect 442604 653880 442728 653980
rect 442828 653880 442952 653980
rect 443052 653880 443176 653980
rect 443276 653880 443400 653980
rect 443500 653880 443624 653980
rect 443724 653880 443848 653980
rect 443948 653880 444072 653980
rect 444172 653880 444296 653980
rect 444396 653880 444520 653980
rect 444620 653880 444744 653980
rect 444844 653880 444968 653980
rect 445068 653880 445192 653980
rect 445292 653880 445416 653980
rect 445516 653880 445540 653980
rect 438880 653846 445540 653880
rect 449350 654876 456010 654906
rect 449350 654776 449390 654876
rect 449490 654776 449614 654876
rect 449714 654776 449838 654876
rect 449938 654776 450062 654876
rect 450162 654776 450286 654876
rect 450386 654776 450510 654876
rect 450610 654776 450734 654876
rect 450834 654776 450958 654876
rect 451058 654776 451182 654876
rect 451282 654776 451406 654876
rect 451506 654776 451630 654876
rect 451730 654776 451854 654876
rect 451954 654776 452078 654876
rect 452178 654776 452302 654876
rect 452402 654776 452526 654876
rect 452626 654776 452750 654876
rect 452850 654776 452974 654876
rect 453074 654776 453198 654876
rect 453298 654776 453422 654876
rect 453522 654776 453646 654876
rect 453746 654776 453870 654876
rect 453970 654776 454094 654876
rect 454194 654776 454318 654876
rect 454418 654776 454542 654876
rect 454642 654776 454766 654876
rect 454866 654776 454990 654876
rect 455090 654776 455214 654876
rect 455314 654776 455438 654876
rect 455538 654776 455662 654876
rect 455762 654776 455886 654876
rect 455986 654776 456010 654876
rect 449350 654652 456010 654776
rect 449350 654552 449390 654652
rect 449490 654552 449614 654652
rect 449714 654552 449838 654652
rect 449938 654552 450062 654652
rect 450162 654552 450286 654652
rect 450386 654552 450510 654652
rect 450610 654552 450734 654652
rect 450834 654552 450958 654652
rect 451058 654552 451182 654652
rect 451282 654552 451406 654652
rect 451506 654552 451630 654652
rect 451730 654552 451854 654652
rect 451954 654552 452078 654652
rect 452178 654552 452302 654652
rect 452402 654552 452526 654652
rect 452626 654552 452750 654652
rect 452850 654552 452974 654652
rect 453074 654552 453198 654652
rect 453298 654552 453422 654652
rect 453522 654552 453646 654652
rect 453746 654552 453870 654652
rect 453970 654552 454094 654652
rect 454194 654552 454318 654652
rect 454418 654552 454542 654652
rect 454642 654552 454766 654652
rect 454866 654552 454990 654652
rect 455090 654552 455214 654652
rect 455314 654552 455438 654652
rect 455538 654552 455662 654652
rect 455762 654552 455886 654652
rect 455986 654552 456010 654652
rect 449350 654428 456010 654552
rect 449350 654328 449390 654428
rect 449490 654328 449614 654428
rect 449714 654328 449838 654428
rect 449938 654328 450062 654428
rect 450162 654328 450286 654428
rect 450386 654328 450510 654428
rect 450610 654328 450734 654428
rect 450834 654328 450958 654428
rect 451058 654328 451182 654428
rect 451282 654328 451406 654428
rect 451506 654328 451630 654428
rect 451730 654328 451854 654428
rect 451954 654328 452078 654428
rect 452178 654328 452302 654428
rect 452402 654328 452526 654428
rect 452626 654328 452750 654428
rect 452850 654328 452974 654428
rect 453074 654328 453198 654428
rect 453298 654328 453422 654428
rect 453522 654328 453646 654428
rect 453746 654328 453870 654428
rect 453970 654328 454094 654428
rect 454194 654328 454318 654428
rect 454418 654328 454542 654428
rect 454642 654328 454766 654428
rect 454866 654328 454990 654428
rect 455090 654328 455214 654428
rect 455314 654328 455438 654428
rect 455538 654328 455662 654428
rect 455762 654328 455886 654428
rect 455986 654328 456010 654428
rect 449350 654204 456010 654328
rect 449350 654104 449390 654204
rect 449490 654104 449614 654204
rect 449714 654104 449838 654204
rect 449938 654104 450062 654204
rect 450162 654104 450286 654204
rect 450386 654104 450510 654204
rect 450610 654104 450734 654204
rect 450834 654104 450958 654204
rect 451058 654104 451182 654204
rect 451282 654104 451406 654204
rect 451506 654104 451630 654204
rect 451730 654104 451854 654204
rect 451954 654104 452078 654204
rect 452178 654104 452302 654204
rect 452402 654104 452526 654204
rect 452626 654104 452750 654204
rect 452850 654104 452974 654204
rect 453074 654104 453198 654204
rect 453298 654104 453422 654204
rect 453522 654104 453646 654204
rect 453746 654104 453870 654204
rect 453970 654104 454094 654204
rect 454194 654104 454318 654204
rect 454418 654104 454542 654204
rect 454642 654104 454766 654204
rect 454866 654104 454990 654204
rect 455090 654104 455214 654204
rect 455314 654104 455438 654204
rect 455538 654104 455662 654204
rect 455762 654104 455886 654204
rect 455986 654104 456010 654204
rect 449350 653980 456010 654104
rect 449350 653880 449390 653980
rect 449490 653880 449614 653980
rect 449714 653880 449838 653980
rect 449938 653880 450062 653980
rect 450162 653880 450286 653980
rect 450386 653880 450510 653980
rect 450610 653880 450734 653980
rect 450834 653880 450958 653980
rect 451058 653880 451182 653980
rect 451282 653880 451406 653980
rect 451506 653880 451630 653980
rect 451730 653880 451854 653980
rect 451954 653880 452078 653980
rect 452178 653880 452302 653980
rect 452402 653880 452526 653980
rect 452626 653880 452750 653980
rect 452850 653880 452974 653980
rect 453074 653880 453198 653980
rect 453298 653880 453422 653980
rect 453522 653880 453646 653980
rect 453746 653880 453870 653980
rect 453970 653880 454094 653980
rect 454194 653880 454318 653980
rect 454418 653880 454542 653980
rect 454642 653880 454766 653980
rect 454866 653880 454990 653980
rect 455090 653880 455214 653980
rect 455314 653880 455438 653980
rect 455538 653880 455662 653980
rect 455762 653880 455886 653980
rect 455986 653880 456010 653980
rect 449350 653846 456010 653880
rect 475620 654896 482280 654926
rect 475620 654796 475660 654896
rect 475760 654796 475884 654896
rect 475984 654796 476108 654896
rect 476208 654796 476332 654896
rect 476432 654796 476556 654896
rect 476656 654796 476780 654896
rect 476880 654796 477004 654896
rect 477104 654796 477228 654896
rect 477328 654796 477452 654896
rect 477552 654796 477676 654896
rect 477776 654796 477900 654896
rect 478000 654796 478124 654896
rect 478224 654796 478348 654896
rect 478448 654796 478572 654896
rect 478672 654796 478796 654896
rect 478896 654796 479020 654896
rect 479120 654796 479244 654896
rect 479344 654796 479468 654896
rect 479568 654796 479692 654896
rect 479792 654796 479916 654896
rect 480016 654796 480140 654896
rect 480240 654796 480364 654896
rect 480464 654796 480588 654896
rect 480688 654796 480812 654896
rect 480912 654796 481036 654896
rect 481136 654796 481260 654896
rect 481360 654796 481484 654896
rect 481584 654796 481708 654896
rect 481808 654796 481932 654896
rect 482032 654796 482156 654896
rect 482256 654796 482280 654896
rect 475620 654672 482280 654796
rect 475620 654572 475660 654672
rect 475760 654572 475884 654672
rect 475984 654572 476108 654672
rect 476208 654572 476332 654672
rect 476432 654572 476556 654672
rect 476656 654572 476780 654672
rect 476880 654572 477004 654672
rect 477104 654572 477228 654672
rect 477328 654572 477452 654672
rect 477552 654572 477676 654672
rect 477776 654572 477900 654672
rect 478000 654572 478124 654672
rect 478224 654572 478348 654672
rect 478448 654572 478572 654672
rect 478672 654572 478796 654672
rect 478896 654572 479020 654672
rect 479120 654572 479244 654672
rect 479344 654572 479468 654672
rect 479568 654572 479692 654672
rect 479792 654572 479916 654672
rect 480016 654572 480140 654672
rect 480240 654572 480364 654672
rect 480464 654572 480588 654672
rect 480688 654572 480812 654672
rect 480912 654572 481036 654672
rect 481136 654572 481260 654672
rect 481360 654572 481484 654672
rect 481584 654572 481708 654672
rect 481808 654572 481932 654672
rect 482032 654572 482156 654672
rect 482256 654572 482280 654672
rect 475620 654448 482280 654572
rect 475620 654348 475660 654448
rect 475760 654348 475884 654448
rect 475984 654348 476108 654448
rect 476208 654348 476332 654448
rect 476432 654348 476556 654448
rect 476656 654348 476780 654448
rect 476880 654348 477004 654448
rect 477104 654348 477228 654448
rect 477328 654348 477452 654448
rect 477552 654348 477676 654448
rect 477776 654348 477900 654448
rect 478000 654348 478124 654448
rect 478224 654348 478348 654448
rect 478448 654348 478572 654448
rect 478672 654348 478796 654448
rect 478896 654348 479020 654448
rect 479120 654348 479244 654448
rect 479344 654348 479468 654448
rect 479568 654348 479692 654448
rect 479792 654348 479916 654448
rect 480016 654348 480140 654448
rect 480240 654348 480364 654448
rect 480464 654348 480588 654448
rect 480688 654348 480812 654448
rect 480912 654348 481036 654448
rect 481136 654348 481260 654448
rect 481360 654348 481484 654448
rect 481584 654348 481708 654448
rect 481808 654348 481932 654448
rect 482032 654348 482156 654448
rect 482256 654348 482280 654448
rect 475620 654224 482280 654348
rect 475620 654124 475660 654224
rect 475760 654124 475884 654224
rect 475984 654124 476108 654224
rect 476208 654124 476332 654224
rect 476432 654124 476556 654224
rect 476656 654124 476780 654224
rect 476880 654124 477004 654224
rect 477104 654124 477228 654224
rect 477328 654124 477452 654224
rect 477552 654124 477676 654224
rect 477776 654124 477900 654224
rect 478000 654124 478124 654224
rect 478224 654124 478348 654224
rect 478448 654124 478572 654224
rect 478672 654124 478796 654224
rect 478896 654124 479020 654224
rect 479120 654124 479244 654224
rect 479344 654124 479468 654224
rect 479568 654124 479692 654224
rect 479792 654124 479916 654224
rect 480016 654124 480140 654224
rect 480240 654124 480364 654224
rect 480464 654124 480588 654224
rect 480688 654124 480812 654224
rect 480912 654124 481036 654224
rect 481136 654124 481260 654224
rect 481360 654124 481484 654224
rect 481584 654124 481708 654224
rect 481808 654124 481932 654224
rect 482032 654124 482156 654224
rect 482256 654124 482280 654224
rect 475620 654000 482280 654124
rect 475620 653900 475660 654000
rect 475760 653900 475884 654000
rect 475984 653900 476108 654000
rect 476208 653900 476332 654000
rect 476432 653900 476556 654000
rect 476656 653900 476780 654000
rect 476880 653900 477004 654000
rect 477104 653900 477228 654000
rect 477328 653900 477452 654000
rect 477552 653900 477676 654000
rect 477776 653900 477900 654000
rect 478000 653900 478124 654000
rect 478224 653900 478348 654000
rect 478448 653900 478572 654000
rect 478672 653900 478796 654000
rect 478896 653900 479020 654000
rect 479120 653900 479244 654000
rect 479344 653900 479468 654000
rect 479568 653900 479692 654000
rect 479792 653900 479916 654000
rect 480016 653900 480140 654000
rect 480240 653900 480364 654000
rect 480464 653900 480588 654000
rect 480688 653900 480812 654000
rect 480912 653900 481036 654000
rect 481136 653900 481260 654000
rect 481360 653900 481484 654000
rect 481584 653900 481708 654000
rect 481808 653900 481932 654000
rect 482032 653900 482156 654000
rect 482256 653900 482280 654000
rect 475620 653866 482280 653900
rect 440696 652754 451952 652760
rect 440696 651928 440702 652754
rect 451946 651928 451952 652754
rect 440696 651922 451952 651928
rect 463962 651214 466156 651220
rect 463962 650656 463968 651214
rect 464526 650656 465592 651214
rect 466150 650656 466156 651214
rect 463962 650650 466156 650656
rect 469508 651214 472706 651220
rect 469508 650656 469682 651214
rect 470240 650656 472136 651214
rect 472694 650656 472706 651214
rect 469508 650650 472706 650656
rect 457406 650414 463702 650420
rect 437864 650178 438924 650202
rect 437864 650078 437894 650178
rect 437994 650078 438118 650178
rect 438218 650078 438342 650178
rect 438442 650078 438566 650178
rect 438666 650078 438790 650178
rect 438890 650078 438924 650178
rect 437864 649954 438924 650078
rect 437864 649854 437894 649954
rect 437994 649854 438118 649954
rect 438218 649854 438342 649954
rect 438442 649854 438566 649954
rect 438666 649854 438790 649954
rect 438890 649854 438924 649954
rect 437864 649730 438924 649854
rect 457406 649856 457412 650414
rect 457970 649856 463138 650414
rect 463696 649856 463702 650414
rect 457406 649850 463702 649856
rect 466282 650414 469428 650420
rect 466282 649856 466410 650414
rect 466968 649856 468864 650414
rect 469422 649856 469428 650414
rect 466282 649850 469428 649856
rect 471198 650414 474336 650420
rect 471198 649856 471318 650414
rect 471876 649856 473772 650414
rect 474330 649856 474336 650414
rect 471198 649850 474336 649856
rect 482144 650178 483204 650202
rect 482144 650078 482174 650178
rect 482274 650078 482398 650178
rect 482498 650078 482622 650178
rect 482722 650078 482846 650178
rect 482946 650078 483070 650178
rect 483170 650078 483204 650178
rect 482144 649954 483204 650078
rect 482144 649854 482174 649954
rect 482274 649854 482398 649954
rect 482498 649854 482622 649954
rect 482722 649854 482846 649954
rect 482946 649854 483070 649954
rect 483170 649854 483204 649954
rect 437864 649630 437894 649730
rect 437994 649630 438118 649730
rect 438218 649630 438342 649730
rect 438442 649630 438566 649730
rect 438666 649630 438790 649730
rect 438890 649630 438924 649730
rect 482144 649730 483204 649854
rect 457406 649676 457976 649682
rect 437864 649506 438924 649630
rect 437864 649406 437894 649506
rect 437994 649406 438118 649506
rect 438218 649406 438342 649506
rect 438442 649406 438566 649506
rect 438666 649406 438790 649506
rect 438890 649406 438924 649506
rect 437864 649282 438924 649406
rect 437864 649182 437894 649282
rect 437994 649182 438118 649282
rect 438218 649182 438342 649282
rect 438442 649182 438566 649282
rect 438666 649182 438790 649282
rect 438890 649182 438924 649282
rect 456592 649664 457154 649670
rect 456592 649267 456604 649664
rect 457142 649267 457154 649664
rect 456592 649261 457154 649267
rect 457406 649256 457412 649676
rect 457970 649256 457976 649676
rect 457406 649250 457976 649256
rect 458224 649676 458794 649682
rect 458224 649256 458230 649676
rect 458788 649256 458794 649676
rect 459046 649664 459608 649670
rect 459046 649267 459058 649664
rect 459596 649267 459608 649664
rect 482144 649630 482174 649730
rect 482274 649630 482398 649730
rect 482498 649630 482622 649730
rect 482722 649630 482846 649730
rect 482946 649630 483070 649730
rect 483170 649630 483204 649730
rect 462314 649614 462884 649620
rect 459046 649261 459608 649267
rect 461500 649602 462062 649608
rect 458224 649250 458794 649256
rect 461500 649205 461512 649602
rect 462050 649205 462062 649602
rect 461500 649199 462062 649205
rect 462314 649194 462320 649614
rect 462878 649194 462884 649614
rect 462314 649188 462884 649194
rect 463132 649614 463702 649620
rect 463132 649194 463138 649614
rect 463696 649194 463702 649614
rect 463132 649188 463702 649194
rect 463950 649614 464520 649620
rect 463950 649194 463956 649614
rect 464514 649194 464520 649614
rect 463950 649188 464520 649194
rect 464768 649614 465338 649620
rect 464768 649194 464774 649614
rect 465332 649194 465338 649614
rect 464768 649188 465338 649194
rect 465586 649614 466156 649620
rect 465586 649194 465592 649614
rect 466150 649194 466156 649614
rect 465586 649188 466156 649194
rect 466404 649614 466974 649620
rect 466404 649194 466410 649614
rect 466968 649194 466974 649614
rect 466404 649188 466974 649194
rect 467222 649614 467792 649620
rect 467222 649194 467228 649614
rect 467786 649194 467792 649614
rect 467222 649188 467792 649194
rect 468040 649614 468610 649620
rect 468040 649194 468046 649614
rect 468604 649194 468610 649614
rect 468040 649188 468610 649194
rect 468858 649614 469428 649620
rect 468858 649194 468864 649614
rect 469422 649194 469428 649614
rect 468858 649188 469428 649194
rect 469676 649614 470246 649620
rect 469676 649194 469682 649614
rect 470240 649194 470246 649614
rect 469676 649188 470246 649194
rect 470494 649614 471064 649620
rect 470494 649194 470500 649614
rect 471058 649194 471064 649614
rect 470494 649188 471064 649194
rect 471312 649614 471882 649620
rect 471312 649194 471318 649614
rect 471876 649194 471882 649614
rect 471312 649188 471882 649194
rect 472130 649614 472700 649620
rect 472130 649194 472136 649614
rect 472694 649194 472700 649614
rect 472130 649188 472700 649194
rect 472948 649614 473518 649620
rect 472948 649194 472954 649614
rect 473512 649194 473518 649614
rect 472948 649188 473518 649194
rect 473766 649614 474336 649620
rect 473766 649194 473772 649614
rect 474330 649194 474336 649614
rect 474588 649602 475150 649608
rect 474588 649205 474600 649602
rect 475138 649205 475150 649602
rect 474588 649199 475150 649205
rect 482144 649506 483204 649630
rect 482144 649406 482174 649506
rect 482274 649406 482398 649506
rect 482498 649406 482622 649506
rect 482722 649406 482846 649506
rect 482946 649406 483070 649506
rect 483170 649406 483204 649506
rect 482144 649282 483204 649406
rect 473766 649188 474336 649194
rect 437864 649058 438924 649182
rect 437864 648958 437894 649058
rect 437994 648958 438118 649058
rect 438218 648958 438342 649058
rect 438442 648958 438566 649058
rect 438666 648958 438790 649058
rect 438890 648958 438924 649058
rect 482144 649182 482174 649282
rect 482274 649182 482398 649282
rect 482498 649182 482622 649282
rect 482722 649182 482846 649282
rect 482946 649182 483070 649282
rect 483170 649182 483204 649282
rect 482144 649058 483204 649182
rect 482144 648958 482174 649058
rect 482274 648958 482398 649058
rect 482498 648958 482622 649058
rect 482722 648958 482846 649058
rect 482946 648958 483070 649058
rect 483170 648958 483204 649058
rect 437864 648834 438924 648958
rect 437864 648734 437894 648834
rect 437994 648734 438118 648834
rect 438218 648734 438342 648834
rect 438442 648734 438566 648834
rect 438666 648734 438790 648834
rect 438890 648734 438924 648834
rect 437864 648610 438924 648734
rect 437864 648510 437894 648610
rect 437994 648510 438118 648610
rect 438218 648510 438342 648610
rect 438442 648510 438566 648610
rect 438666 648510 438790 648610
rect 438890 648510 438924 648610
rect 437864 648386 438924 648510
rect 458222 648952 462884 648958
rect 458222 648460 458230 648952
rect 458788 648460 462320 648952
rect 458222 648394 462320 648460
rect 462878 648394 462884 648952
rect 458222 648388 462884 648394
rect 464768 648952 467792 648958
rect 464768 648394 464774 648952
rect 465332 648394 467228 648952
rect 467786 648394 467792 648952
rect 464768 648388 467792 648394
rect 470494 648952 473518 648958
rect 470494 648394 470500 648952
rect 471058 648394 472954 648952
rect 473512 648394 473518 648952
rect 470494 648388 473518 648394
rect 482144 648834 483204 648958
rect 482144 648734 482174 648834
rect 482274 648734 482398 648834
rect 482498 648734 482622 648834
rect 482722 648734 482846 648834
rect 482946 648734 483070 648834
rect 483170 648734 483204 648834
rect 482144 648610 483204 648734
rect 482144 648510 482174 648610
rect 482274 648510 482398 648610
rect 482498 648510 482622 648610
rect 482722 648510 482846 648610
rect 482946 648510 483070 648610
rect 483170 648510 483204 648610
rect 437864 648286 437894 648386
rect 437994 648286 438118 648386
rect 438218 648286 438342 648386
rect 438442 648286 438566 648386
rect 438666 648286 438790 648386
rect 438890 648286 438924 648386
rect 437864 648162 438924 648286
rect 482144 648386 483204 648510
rect 482144 648286 482174 648386
rect 482274 648286 482398 648386
rect 482498 648286 482622 648386
rect 482722 648286 482846 648386
rect 482946 648286 483070 648386
rect 483170 648286 483204 648386
rect 437864 648062 437894 648162
rect 437994 648062 438118 648162
rect 438218 648062 438342 648162
rect 438442 648062 438566 648162
rect 438666 648062 438790 648162
rect 438890 648062 438924 648162
rect 437864 647938 438924 648062
rect 437864 647838 437894 647938
rect 437994 647838 438118 647938
rect 438218 647838 438342 647938
rect 438442 647838 438566 647938
rect 438666 647838 438790 647938
rect 438890 647838 438924 647938
rect 453320 648278 453882 648284
rect 453320 647881 453332 648278
rect 453870 647881 453882 648278
rect 453320 647875 453882 647881
rect 454138 648278 454700 648284
rect 454138 647881 454150 648278
rect 454688 647881 454700 648278
rect 454138 647875 454700 647881
rect 454956 648278 455518 648284
rect 454956 647881 454968 648278
rect 455506 647881 455518 648278
rect 454956 647875 455518 647881
rect 482144 648162 483204 648286
rect 482144 648062 482174 648162
rect 482274 648062 482398 648162
rect 482498 648062 482622 648162
rect 482722 648062 482846 648162
rect 482946 648062 483070 648162
rect 483170 648062 483204 648162
rect 482144 647938 483204 648062
rect 437864 647714 438924 647838
rect 437864 647614 437894 647714
rect 437994 647614 438118 647714
rect 438218 647614 438342 647714
rect 438442 647614 438566 647714
rect 438666 647614 438790 647714
rect 438890 647614 438924 647714
rect 437864 647490 438924 647614
rect 437864 647390 437894 647490
rect 437994 647390 438118 647490
rect 438218 647390 438342 647490
rect 438442 647390 438566 647490
rect 438666 647390 438790 647490
rect 438890 647390 438924 647490
rect 437864 647266 438924 647390
rect 437864 647166 437894 647266
rect 437994 647166 438118 647266
rect 438218 647166 438342 647266
rect 438442 647166 438566 647266
rect 438666 647166 438790 647266
rect 438890 647166 438924 647266
rect 437864 647042 438924 647166
rect 437864 646942 437894 647042
rect 437994 646942 438118 647042
rect 438218 646942 438342 647042
rect 438442 646942 438566 647042
rect 438666 646942 438790 647042
rect 438890 646942 438924 647042
rect 437864 646818 438924 646942
rect 437864 646718 437894 646818
rect 437994 646718 438118 646818
rect 438218 646718 438342 646818
rect 438442 646718 438566 646818
rect 438666 646718 438790 646818
rect 438890 646718 438924 646818
rect 437864 646594 438924 646718
rect 437864 646494 437894 646594
rect 437994 646494 438118 646594
rect 438218 646494 438342 646594
rect 438442 646494 438566 646594
rect 438666 646494 438790 646594
rect 438890 646494 438924 646594
rect 437864 646370 438924 646494
rect 437864 646270 437894 646370
rect 437994 646270 438118 646370
rect 438218 646270 438342 646370
rect 438442 646270 438566 646370
rect 438666 646270 438790 646370
rect 438890 646270 438924 646370
rect 437864 646146 438924 646270
rect 437864 646046 437894 646146
rect 437994 646046 438118 646146
rect 438218 646046 438342 646146
rect 438442 646046 438566 646146
rect 438666 646046 438790 646146
rect 438890 646046 438924 646146
rect 437864 645922 438924 646046
rect 437864 645822 437894 645922
rect 437994 645822 438118 645922
rect 438218 645822 438342 645922
rect 438442 645822 438566 645922
rect 438666 645822 438790 645922
rect 438890 645822 438924 645922
rect 437864 645698 438924 645822
rect 437864 645598 437894 645698
rect 437994 645598 438118 645698
rect 438218 645598 438342 645698
rect 438442 645598 438566 645698
rect 438666 645598 438790 645698
rect 438890 645598 438924 645698
rect 437864 645474 438924 645598
rect 437864 645374 437894 645474
rect 437994 645374 438118 645474
rect 438218 645374 438342 645474
rect 438442 645374 438566 645474
rect 438666 645374 438790 645474
rect 438890 645374 438924 645474
rect 437864 645250 438924 645374
rect 437864 645150 437894 645250
rect 437994 645150 438118 645250
rect 438218 645150 438342 645250
rect 438442 645150 438566 645250
rect 438666 645150 438790 645250
rect 438890 645150 438924 645250
rect 437864 645026 438924 645150
rect 437864 644926 437894 645026
rect 437994 644926 438118 645026
rect 438218 644926 438342 645026
rect 438442 644926 438566 645026
rect 438666 644926 438790 645026
rect 438890 644926 438924 645026
rect 482144 647838 482174 647938
rect 482274 647838 482398 647938
rect 482498 647838 482622 647938
rect 482722 647838 482846 647938
rect 482946 647838 483070 647938
rect 483170 647838 483204 647938
rect 482144 647714 483204 647838
rect 482144 647614 482174 647714
rect 482274 647614 482398 647714
rect 482498 647614 482622 647714
rect 482722 647614 482846 647714
rect 482946 647614 483070 647714
rect 483170 647614 483204 647714
rect 482144 647490 483204 647614
rect 482144 647390 482174 647490
rect 482274 647390 482398 647490
rect 482498 647390 482622 647490
rect 482722 647390 482846 647490
rect 482946 647390 483070 647490
rect 483170 647390 483204 647490
rect 482144 647266 483204 647390
rect 482144 647166 482174 647266
rect 482274 647166 482398 647266
rect 482498 647166 482622 647266
rect 482722 647166 482846 647266
rect 482946 647166 483070 647266
rect 483170 647166 483204 647266
rect 482144 647042 483204 647166
rect 482144 646942 482174 647042
rect 482274 646942 482398 647042
rect 482498 646942 482622 647042
rect 482722 646942 482846 647042
rect 482946 646942 483070 647042
rect 483170 646942 483204 647042
rect 482144 646818 483204 646942
rect 482144 646718 482174 646818
rect 482274 646718 482398 646818
rect 482498 646718 482622 646818
rect 482722 646718 482846 646818
rect 482946 646718 483070 646818
rect 483170 646718 483204 646818
rect 482144 646594 483204 646718
rect 482144 646494 482174 646594
rect 482274 646494 482398 646594
rect 482498 646494 482622 646594
rect 482722 646494 482846 646594
rect 482946 646494 483070 646594
rect 483170 646494 483204 646594
rect 482144 646370 483204 646494
rect 482144 646270 482174 646370
rect 482274 646270 482398 646370
rect 482498 646270 482622 646370
rect 482722 646270 482846 646370
rect 482946 646270 483070 646370
rect 483170 646270 483204 646370
rect 482144 646146 483204 646270
rect 482144 646046 482174 646146
rect 482274 646046 482398 646146
rect 482498 646046 482622 646146
rect 482722 646046 482846 646146
rect 482946 646046 483070 646146
rect 483170 646046 483204 646146
rect 482144 645922 483204 646046
rect 482144 645822 482174 645922
rect 482274 645822 482398 645922
rect 482498 645822 482622 645922
rect 482722 645822 482846 645922
rect 482946 645822 483070 645922
rect 483170 645822 483204 645922
rect 482144 645698 483204 645822
rect 482144 645598 482174 645698
rect 482274 645598 482398 645698
rect 482498 645598 482622 645698
rect 482722 645598 482846 645698
rect 482946 645598 483070 645698
rect 483170 645598 483204 645698
rect 482144 645474 483204 645598
rect 482144 645374 482174 645474
rect 482274 645374 482398 645474
rect 482498 645374 482622 645474
rect 482722 645374 482846 645474
rect 482946 645374 483070 645474
rect 483170 645374 483204 645474
rect 482144 645250 483204 645374
rect 482144 645150 482174 645250
rect 482274 645150 482398 645250
rect 482498 645150 482622 645250
rect 482722 645150 482846 645250
rect 482946 645150 483070 645250
rect 483170 645150 483204 645250
rect 482144 645026 483204 645150
rect 437864 644802 438924 644926
rect 437864 644702 437894 644802
rect 437994 644702 438118 644802
rect 438218 644702 438342 644802
rect 438442 644702 438566 644802
rect 438666 644702 438790 644802
rect 438890 644702 438924 644802
rect 437864 644578 438924 644702
rect 437864 644478 437894 644578
rect 437994 644478 438118 644578
rect 438218 644478 438342 644578
rect 438442 644478 438566 644578
rect 438666 644478 438790 644578
rect 438890 644478 438924 644578
rect 455766 644933 461262 644950
rect 455766 644922 456604 644933
rect 437864 644354 438924 644478
rect 437864 644254 437894 644354
rect 437994 644254 438118 644354
rect 438218 644254 438342 644354
rect 438442 644254 438566 644354
rect 438666 644254 438790 644354
rect 438890 644254 438924 644354
rect 437864 644130 438924 644254
rect 437864 644030 437894 644130
rect 437994 644030 438118 644130
rect 438218 644030 438342 644130
rect 438442 644030 438566 644130
rect 438666 644030 438790 644130
rect 438890 644030 438924 644130
rect 453320 644523 453882 644529
rect 453320 644126 453332 644523
rect 453870 644126 453882 644523
rect 453320 644120 453882 644126
rect 454134 644523 454704 644540
rect 454134 644126 454150 644523
rect 454688 644126 454704 644523
rect 437864 643906 438924 644030
rect 437864 643806 437894 643906
rect 437994 643806 438118 643906
rect 438218 643806 438342 643906
rect 438442 643806 438566 643906
rect 438666 643806 438790 643906
rect 438890 643806 438924 643906
rect 437864 643682 438924 643806
rect 437864 643582 437894 643682
rect 437994 643582 438118 643682
rect 438218 643582 438342 643682
rect 438442 643582 438566 643682
rect 438666 643582 438790 643682
rect 438890 643582 438924 643682
rect 437864 643542 438924 643582
rect 454134 643684 454704 644126
rect 454956 644523 455518 644529
rect 454956 644126 454968 644523
rect 455506 644126 455518 644523
rect 454956 644120 455518 644126
rect 455766 643856 455788 644922
rect 456282 644536 456604 644922
rect 457142 644536 457422 644933
rect 457960 644536 458240 644933
rect 458778 644536 459058 644933
rect 459596 644920 461262 644933
rect 459596 644536 460740 644920
rect 456282 643868 460740 644536
rect 461252 643868 461262 644920
rect 482144 644926 482174 645026
rect 482274 644926 482398 645026
rect 482498 644926 482622 645026
rect 482722 644926 482846 645026
rect 482946 644926 483070 645026
rect 483170 644926 483204 645026
rect 482144 644802 483204 644926
rect 482144 644702 482174 644802
rect 482274 644702 482398 644802
rect 482498 644702 482622 644802
rect 482722 644702 482846 644802
rect 482946 644702 483070 644802
rect 483170 644702 483204 644802
rect 482144 644578 483204 644702
rect 463132 644478 466974 644484
rect 463132 643920 463138 644478
rect 463696 643920 466410 644478
rect 466968 643920 466974 644478
rect 463132 643914 466974 643920
rect 468864 644478 471882 644484
rect 469422 643920 471318 644478
rect 471876 643920 471882 644478
rect 468864 643914 471882 643920
rect 482144 644478 482174 644578
rect 482274 644478 482398 644578
rect 482498 644478 482622 644578
rect 482722 644478 482846 644578
rect 482946 644478 483070 644578
rect 483170 644478 483204 644578
rect 482144 644354 483204 644478
rect 482144 644254 482174 644354
rect 482274 644254 482398 644354
rect 482498 644254 482622 644354
rect 482722 644254 482846 644354
rect 482946 644254 483070 644354
rect 483170 644254 483204 644354
rect 482144 644130 483204 644254
rect 482144 644030 482174 644130
rect 482274 644030 482398 644130
rect 482498 644030 482622 644130
rect 482722 644030 482846 644130
rect 482946 644030 483070 644130
rect 483170 644030 483204 644130
rect 456282 643856 461262 643868
rect 455766 643814 461262 643856
rect 482144 643906 483204 644030
rect 482144 643806 482174 643906
rect 482274 643806 482398 643906
rect 482498 643806 482622 643906
rect 482722 643806 482846 643906
rect 482946 643806 483070 643906
rect 483170 643806 483204 643906
rect 454134 643678 464520 643684
rect 454134 643120 463956 643678
rect 464514 643120 464520 643678
rect 454134 643114 464520 643120
rect 465586 643678 470246 643684
rect 465586 643120 465592 643678
rect 466150 643120 469682 643678
rect 470240 643120 470246 643678
rect 482144 643682 483204 643806
rect 482144 643582 482174 643682
rect 482274 643582 482398 643682
rect 482498 643582 482622 643682
rect 482722 643582 482846 643682
rect 482946 643582 483070 643682
rect 483170 643582 483204 643682
rect 482144 643542 483204 643582
rect 465586 643114 470246 643120
rect 462314 642878 462884 642884
rect 461500 642867 462062 642873
rect 461500 642470 461512 642867
rect 462050 642470 462062 642867
rect 461500 642464 462062 642470
rect 462314 642458 462320 642878
rect 462878 642458 462884 642878
rect 462314 642452 462884 642458
rect 463132 642878 463702 642884
rect 463132 642458 463138 642878
rect 463696 642458 463702 642878
rect 463132 642452 463702 642458
rect 463950 642878 464520 642884
rect 463950 642458 463956 642878
rect 464514 642458 464520 642878
rect 463950 642452 464520 642458
rect 464768 642878 465338 642884
rect 464768 642458 464774 642878
rect 465332 642458 465338 642878
rect 464768 642452 465338 642458
rect 465586 642878 466156 642884
rect 465586 642458 465592 642878
rect 466150 642458 466156 642878
rect 465586 642452 466156 642458
rect 466404 642878 466974 642884
rect 466404 642458 466410 642878
rect 466968 642458 466974 642878
rect 466404 642452 466974 642458
rect 467222 642878 467792 642884
rect 467222 642458 467228 642878
rect 467786 642458 467792 642878
rect 467222 642452 467792 642458
rect 467962 642878 468666 642884
rect 467962 642846 468046 642878
rect 467962 642328 467968 642846
rect 468604 642846 468666 642878
rect 468660 642328 468666 642846
rect 468858 642878 469428 642884
rect 468858 642458 468864 642878
rect 469422 642458 469428 642878
rect 468858 642452 469428 642458
rect 469676 642878 470246 642884
rect 469676 642458 469682 642878
rect 470240 642458 470246 642878
rect 469676 642452 470246 642458
rect 470494 642878 471064 642884
rect 470494 642458 470500 642878
rect 471058 642458 471064 642878
rect 470494 642452 471064 642458
rect 471312 642878 471882 642884
rect 471312 642458 471318 642878
rect 471876 642458 471882 642878
rect 471312 642452 471882 642458
rect 472052 642878 472756 642884
rect 462314 642216 465338 642222
rect 462314 641658 462320 642216
rect 462878 641658 464774 642216
rect 465332 641658 465338 642216
rect 462314 641652 465338 641658
rect 467222 642216 471064 642222
rect 467222 641658 467228 642216
rect 467786 641658 470500 642216
rect 471058 641658 471064 642216
rect 467222 641652 471064 641658
rect 472052 642186 472058 642878
rect 472750 642186 472756 642878
rect 472052 641188 472756 642186
rect 459358 641050 472756 641188
rect 459358 640850 459444 641050
rect 459644 640850 459878 641050
rect 460078 640850 460312 641050
rect 460512 640850 460746 641050
rect 460946 640850 461180 641050
rect 461380 640850 461614 641050
rect 461814 640850 462048 641050
rect 462248 640850 462482 641050
rect 462682 640850 462916 641050
rect 463116 640850 463350 641050
rect 463550 640850 463784 641050
rect 463984 640850 464184 641050
rect 464384 640850 464584 641050
rect 464784 640850 464984 641050
rect 465184 640850 465384 641050
rect 465584 640850 465784 641050
rect 465984 640850 466184 641050
rect 466384 640850 466584 641050
rect 466784 640850 466984 641050
rect 467184 640850 467384 641050
rect 467584 640850 468984 641050
rect 469184 640850 469384 641050
rect 469584 640850 469784 641050
rect 469984 640850 470184 641050
rect 470384 640850 470584 641050
rect 470784 640850 470984 641050
rect 471184 640850 471384 641050
rect 471584 640850 471784 641050
rect 471984 640850 472184 641050
rect 472384 640850 472756 641050
rect 459358 640616 472756 640850
rect 459358 640416 459444 640616
rect 459644 640416 459878 640616
rect 460078 640416 460312 640616
rect 460512 640416 460746 640616
rect 460946 640416 461180 640616
rect 461380 640416 461614 640616
rect 461814 640416 462048 640616
rect 462248 640416 462482 640616
rect 462682 640416 462916 640616
rect 463116 640416 463350 640616
rect 463550 640416 463784 640616
rect 463984 640496 472756 640616
rect 472870 642878 473574 642884
rect 472870 642186 472876 642878
rect 473568 642186 473574 642878
rect 463984 640416 464058 640496
rect 459358 640182 464058 640416
rect 459358 639982 459444 640182
rect 459644 639982 459878 640182
rect 460078 639982 460312 640182
rect 460512 639982 460746 640182
rect 460946 639982 461180 640182
rect 461380 639982 461614 640182
rect 461814 639982 462048 640182
rect 462248 639982 462482 640182
rect 462682 639982 462916 640182
rect 463116 639982 463350 640182
rect 463550 639982 463784 640182
rect 463984 639982 464058 640182
rect 453858 639548 455858 639590
rect 453858 639098 453864 639548
rect 455852 639098 455858 639548
rect 452340 638792 452472 638798
rect 452340 638378 452346 638792
rect 452466 638378 452472 638792
rect 451884 638086 452016 638372
rect 451884 637794 451890 638086
rect 452010 637794 452016 638086
rect 444348 637076 450836 637088
rect 437864 636778 438922 636788
rect 437864 636678 437894 636778
rect 437994 636678 438118 636778
rect 438218 636678 438342 636778
rect 438442 636678 438566 636778
rect 438666 636678 438790 636778
rect 438890 636678 438922 636778
rect 437864 636554 438922 636678
rect 437864 636454 437894 636554
rect 437994 636454 438118 636554
rect 438218 636454 438342 636554
rect 438442 636454 438566 636554
rect 438666 636454 438790 636554
rect 438890 636454 438922 636554
rect 444348 636732 444360 637076
rect 450824 636732 450836 637076
rect 444348 636540 450836 636732
rect 444348 636520 445084 636540
rect 445072 636506 445084 636520
rect 450460 636520 450836 636540
rect 450460 636506 450472 636520
rect 445072 636500 450472 636506
rect 437864 636330 438922 636454
rect 437864 636230 437894 636330
rect 437994 636230 438118 636330
rect 438218 636230 438342 636330
rect 438442 636230 438566 636330
rect 438666 636230 438790 636330
rect 438890 636230 438922 636330
rect 437864 636106 438922 636230
rect 442994 636386 445040 636398
rect 442994 636366 445000 636386
rect 442994 636296 443016 636366
rect 443076 636296 443088 636366
rect 443148 636296 443160 636366
rect 443220 636296 443232 636366
rect 443292 636296 443304 636366
rect 443364 636296 443376 636366
rect 443436 636296 443448 636366
rect 443508 636296 443520 636366
rect 443580 636296 445000 636366
rect 442994 636272 445000 636296
rect 442994 636202 443016 636272
rect 443076 636202 443088 636272
rect 443148 636202 443160 636272
rect 443220 636202 443232 636272
rect 443292 636202 443304 636272
rect 443364 636202 443376 636272
rect 443436 636202 443448 636272
rect 443508 636202 443520 636272
rect 443580 636202 445000 636272
rect 445034 636202 445040 636386
rect 442994 636190 445040 636202
rect 437864 636006 437894 636106
rect 437994 636006 438118 636106
rect 438218 636006 438342 636106
rect 438442 636006 438566 636106
rect 438666 636006 438790 636106
rect 438890 636006 438922 636106
rect 445072 636082 450472 636088
rect 437864 635882 438922 636006
rect 437864 635782 437894 635882
rect 437994 635782 438118 635882
rect 438218 635782 438342 635882
rect 438442 635782 438566 635882
rect 438666 635782 438790 635882
rect 438890 635782 438922 635882
rect 437864 635658 438922 635782
rect 437864 635558 437894 635658
rect 437994 635558 438118 635658
rect 438218 635558 438342 635658
rect 438442 635558 438566 635658
rect 438666 635558 438790 635658
rect 438890 635558 438922 635658
rect 437864 635434 438922 635558
rect 437864 635334 437894 635434
rect 437994 635334 438118 635434
rect 438218 635334 438342 635434
rect 438442 635334 438566 635434
rect 438666 635334 438790 635434
rect 438890 635334 438922 635434
rect 437864 635210 438922 635334
rect 437864 635110 437894 635210
rect 437994 635110 438118 635210
rect 438218 635110 438342 635210
rect 438442 635110 438566 635210
rect 438666 635110 438790 635210
rect 438890 635110 438922 635210
rect 437864 634986 438922 635110
rect 437864 634886 437894 634986
rect 437994 634886 438118 634986
rect 438218 634886 438342 634986
rect 438442 634886 438566 634986
rect 438666 634886 438790 634986
rect 438890 634886 438922 634986
rect 437864 634762 438922 634886
rect 437864 634662 437894 634762
rect 437994 634662 438118 634762
rect 438218 634662 438342 634762
rect 438442 634662 438566 634762
rect 438666 634662 438790 634762
rect 438890 634662 438922 634762
rect 437864 634538 438922 634662
rect 437864 634438 437894 634538
rect 437994 634438 438118 634538
rect 438218 634438 438342 634538
rect 438442 634438 438566 634538
rect 438666 634438 438790 634538
rect 438890 634438 438922 634538
rect 437864 634314 438922 634438
rect 437864 634214 437894 634314
rect 437994 634214 438118 634314
rect 438218 634214 438342 634314
rect 438442 634214 438566 634314
rect 438666 634214 438790 634314
rect 438890 634214 438922 634314
rect 437864 634090 438922 634214
rect 437864 633990 437894 634090
rect 437994 633990 438118 634090
rect 438218 633990 438342 634090
rect 438442 633990 438566 634090
rect 438666 633990 438790 634090
rect 438890 633990 438922 634090
rect 437864 633866 438922 633990
rect 437864 633766 437894 633866
rect 437994 633766 438118 633866
rect 438218 633766 438342 633866
rect 438442 633766 438566 633866
rect 438666 633766 438790 633866
rect 438890 633766 438922 633866
rect 437864 633642 438922 633766
rect 437864 633542 437894 633642
rect 437994 633542 438118 633642
rect 438218 633542 438342 633642
rect 438442 633542 438566 633642
rect 438666 633542 438790 633642
rect 438890 633542 438922 633642
rect 437864 633418 438922 633542
rect 444354 636048 445084 636082
rect 450460 636048 450830 636082
rect 444354 635726 450830 636048
rect 437864 633318 437894 633418
rect 437994 633318 438118 633418
rect 438218 633318 438342 633418
rect 438442 633318 438566 633418
rect 438666 633318 438790 633418
rect 438890 633318 438922 633418
rect 441330 633408 441406 633420
rect 441330 633356 441342 633408
rect 441394 633356 441406 633408
rect 441330 633344 441406 633356
rect 442246 633408 442322 633420
rect 442246 633356 442258 633408
rect 442310 633356 442322 633408
rect 442246 633344 442322 633356
rect 437864 633194 438922 633318
rect 440578 633292 440786 633298
rect 441024 633292 441256 633304
rect 440578 633258 440590 633292
rect 440774 633258 440786 633292
rect 440578 633252 440786 633258
rect 440888 633258 441048 633292
rect 441232 633258 441256 633292
rect 440888 633220 440932 633258
rect 441024 633240 441256 633258
rect 437864 633094 437894 633194
rect 437994 633094 438118 633194
rect 438218 633094 438342 633194
rect 438442 633094 438566 633194
rect 438666 633094 438790 633194
rect 438890 633094 438922 633194
rect 437864 632970 438922 633094
rect 437864 632870 437894 632970
rect 437994 632870 438118 632970
rect 438218 632870 438342 632970
rect 438442 632870 438566 632970
rect 438666 632870 438790 632970
rect 438890 632870 438922 632970
rect 437864 632746 438922 632870
rect 440430 633208 440476 633220
rect 440430 632832 440436 633208
rect 440470 632832 440476 633208
rect 440430 632820 440476 632832
rect 440888 633208 440934 633220
rect 440888 632832 440894 633208
rect 440928 632832 440934 633208
rect 437864 632646 437894 632746
rect 437994 632646 438118 632746
rect 438218 632646 438342 632746
rect 438442 632646 438566 632746
rect 438666 632646 438790 632746
rect 438890 632646 438922 632746
rect 440888 632690 440934 632832
rect 441346 633208 441392 633344
rect 441494 633292 441702 633298
rect 441494 633258 441506 633292
rect 441690 633258 441702 633292
rect 441494 633252 441702 633258
rect 441952 633292 442160 633298
rect 441952 633258 441964 633292
rect 442148 633258 442160 633292
rect 441952 633252 442160 633258
rect 441346 632832 441352 633208
rect 441386 632832 441392 633208
rect 441346 632820 441392 632832
rect 441804 633208 441850 633220
rect 441804 632832 441810 633208
rect 441844 632832 441850 633208
rect 437864 632522 438922 632646
rect 440878 632684 440942 632690
rect 440878 632632 440884 632684
rect 440936 632632 440942 632684
rect 440878 632626 440942 632632
rect 437864 632422 437894 632522
rect 437994 632422 438118 632522
rect 438218 632422 438342 632522
rect 438442 632422 438566 632522
rect 438666 632422 438790 632522
rect 438890 632422 438922 632522
rect 441804 632484 441850 632832
rect 442262 633208 442308 633344
rect 442388 633292 442620 633304
rect 442868 633292 443076 633298
rect 442388 633258 442422 633292
rect 442606 633258 442766 633292
rect 442388 633240 442620 633258
rect 442262 632832 442268 633208
rect 442302 632832 442308 633208
rect 442262 632820 442308 632832
rect 442720 633208 442766 633258
rect 442868 633258 442880 633292
rect 443064 633258 443076 633292
rect 442868 633252 443076 633258
rect 442720 632832 442726 633208
rect 442760 632832 442766 633208
rect 442720 632696 442766 632832
rect 443178 633208 443224 633220
rect 443178 632832 443184 633208
rect 443218 632832 443224 633208
rect 443178 632820 443224 632832
rect 442712 632690 442776 632696
rect 442712 632638 442718 632690
rect 442770 632638 442776 632690
rect 442712 632632 442776 632638
rect 443318 632690 443524 632696
rect 443318 632632 443324 632690
rect 443518 632632 443524 632690
rect 437864 632298 438922 632422
rect 441796 632478 441860 632484
rect 441796 632426 441802 632478
rect 441854 632426 441860 632478
rect 441796 632420 441860 632426
rect 437864 632198 437894 632298
rect 437994 632198 438118 632298
rect 438218 632198 438342 632298
rect 438442 632198 438566 632298
rect 438666 632198 438790 632298
rect 438890 632198 438922 632298
rect 437864 632074 438922 632198
rect 437864 631974 437894 632074
rect 437994 631974 438118 632074
rect 438218 631974 438342 632074
rect 438442 631974 438566 632074
rect 438666 631974 438790 632074
rect 438890 631974 438922 632074
rect 437864 631850 438922 631974
rect 437864 631750 437894 631850
rect 437994 631750 438118 631850
rect 438218 631750 438342 631850
rect 438442 631750 438566 631850
rect 438666 631750 438790 631850
rect 438890 631750 438922 631850
rect 437864 631626 438922 631750
rect 437864 631526 437894 631626
rect 437994 631526 438118 631626
rect 438218 631526 438342 631626
rect 438442 631526 438566 631626
rect 438666 631526 438790 631626
rect 438890 631526 438922 631626
rect 437864 631402 438922 631526
rect 437864 631302 437894 631402
rect 437994 631302 438118 631402
rect 438218 631302 438342 631402
rect 438442 631302 438566 631402
rect 438666 631302 438790 631402
rect 438890 631302 438922 631402
rect 437864 631178 438922 631302
rect 437864 631078 437894 631178
rect 437994 631078 438118 631178
rect 438218 631078 438342 631178
rect 438442 631078 438566 631178
rect 438666 631078 438790 631178
rect 438890 631078 438922 631178
rect 437864 630954 438922 631078
rect 437864 630854 437894 630954
rect 437994 630854 438118 630954
rect 438218 630854 438342 630954
rect 438442 630854 438566 630954
rect 438666 630854 438790 630954
rect 438890 630854 438922 630954
rect 437864 630730 438922 630854
rect 437864 630630 437894 630730
rect 437994 630630 438118 630730
rect 438218 630630 438342 630730
rect 438442 630630 438566 630730
rect 438666 630630 438790 630730
rect 438890 630630 438922 630730
rect 437864 630506 438922 630630
rect 437864 630406 437894 630506
rect 437994 630406 438118 630506
rect 438218 630406 438342 630506
rect 438442 630406 438566 630506
rect 438666 630406 438790 630506
rect 438890 630406 438922 630506
rect 437864 630282 438922 630406
rect 437864 630182 437894 630282
rect 437994 630182 438118 630282
rect 438218 630182 438342 630282
rect 438442 630182 438566 630282
rect 438666 630182 438790 630282
rect 438890 630182 438922 630282
rect 437864 630162 438922 630182
rect 442982 631830 443114 631842
rect 442982 629488 442998 631830
rect 443098 629488 443114 631830
rect 442982 629240 443114 629488
rect 442982 629136 443008 629240
rect 443060 629136 443114 629240
rect 442982 629126 443114 629136
rect 443318 629046 443524 632632
rect 444354 632318 444562 635726
rect 446664 634674 446848 634694
rect 446664 634620 446684 634674
rect 446828 634620 446848 634674
rect 446092 634534 446276 634554
rect 446092 634480 446112 634534
rect 446256 634480 446276 634534
rect 446092 634420 446276 634480
rect 446664 634420 446848 634620
rect 447808 634674 447992 634694
rect 447808 634620 447828 634674
rect 447972 634620 447992 634674
rect 447236 634534 447420 634554
rect 447236 634480 447256 634534
rect 447400 634480 447420 634534
rect 447236 634420 447420 634480
rect 447808 634420 447992 634620
rect 448952 634674 449136 634694
rect 448952 634620 448972 634674
rect 449116 634620 449136 634674
rect 448380 634534 448564 634554
rect 448380 634480 448400 634534
rect 448544 634480 448564 634534
rect 448380 634420 448564 634480
rect 448952 634420 449136 634620
rect 444808 634414 445864 634420
rect 444808 634380 445520 634414
rect 445704 634380 445864 634414
rect 444808 634374 445864 634380
rect 446080 634414 446288 634420
rect 446080 634380 446092 634414
rect 446276 634380 446288 634414
rect 446080 634374 446288 634380
rect 446652 634414 446860 634420
rect 446652 634380 446664 634414
rect 446848 634380 446860 634414
rect 446652 634374 446860 634380
rect 447224 634414 447432 634420
rect 447224 634380 447236 634414
rect 447420 634380 447432 634414
rect 447224 634374 447432 634380
rect 447796 634414 448004 634420
rect 447796 634380 447808 634414
rect 447992 634380 448004 634414
rect 447796 634374 448004 634380
rect 448368 634414 448576 634420
rect 448368 634380 448380 634414
rect 448564 634380 448576 634414
rect 448368 634374 448576 634380
rect 448940 634414 449148 634420
rect 448940 634380 448952 634414
rect 449136 634380 449148 634414
rect 448940 634374 449148 634380
rect 449364 634414 450420 634420
rect 449364 634380 449524 634414
rect 449708 634380 450420 634414
rect 449364 634374 450420 634380
rect 444808 634346 444922 634374
rect 444798 634330 444930 634346
rect 444798 632732 444814 634330
rect 444914 632732 444930 634330
rect 444798 632714 444930 632732
rect 445360 634330 445406 634374
rect 445360 632554 445366 634330
rect 445400 632554 445406 634330
rect 445360 632542 445406 632554
rect 445818 634330 445864 634374
rect 445818 632554 445824 634330
rect 445858 632554 445864 634330
rect 445818 632542 445864 632554
rect 445932 634330 445978 634342
rect 445932 632554 445938 634330
rect 445972 632554 445978 634330
rect 445932 632542 445978 632554
rect 446390 634330 446436 634342
rect 446390 632554 446396 634330
rect 446430 632554 446436 634330
rect 446390 632542 446436 632554
rect 446504 634330 446550 634342
rect 446504 632554 446510 634330
rect 446544 632554 446550 634330
rect 446504 632542 446550 632554
rect 446962 634330 447008 634342
rect 446962 632554 446968 634330
rect 447002 632554 447008 634330
rect 446962 632542 447008 632554
rect 447076 634330 447122 634342
rect 447076 632554 447082 634330
rect 447116 632554 447122 634330
rect 447076 632542 447122 632554
rect 447534 634330 447580 634342
rect 447534 632554 447540 634330
rect 447574 632554 447580 634330
rect 447534 632542 447580 632554
rect 447648 634330 447694 634342
rect 447648 632554 447654 634330
rect 447688 632554 447694 634330
rect 447648 632542 447694 632554
rect 448106 634330 448152 634342
rect 448106 632554 448112 634330
rect 448146 632554 448152 634330
rect 448106 632542 448152 632554
rect 448220 634330 448266 634342
rect 448220 632554 448226 634330
rect 448260 632554 448266 634330
rect 448220 632542 448266 632554
rect 448678 634330 448724 634342
rect 448678 632554 448684 634330
rect 448718 632554 448724 634330
rect 448678 632542 448724 632554
rect 448792 634330 448838 634342
rect 448792 632554 448798 634330
rect 448832 632554 448838 634330
rect 448792 632542 448838 632554
rect 449250 634330 449296 634342
rect 449250 632554 449256 634330
rect 449290 632554 449296 634330
rect 449250 632542 449296 632554
rect 449364 634330 449410 634374
rect 449364 632554 449370 634330
rect 449404 632554 449410 634330
rect 449364 632542 449410 632554
rect 449822 634330 449868 634374
rect 450306 634346 450420 634374
rect 449822 632554 449828 634330
rect 449862 632554 449868 634330
rect 450298 634330 450430 634346
rect 450298 632732 450314 634330
rect 450414 632732 450430 634330
rect 450298 632714 450430 632732
rect 449822 632542 449868 632554
rect 444354 632064 444480 632318
rect 444532 632064 444562 632318
rect 443634 632011 444138 632018
rect 443634 631977 443794 632011
rect 443978 631977 444138 632011
rect 443634 631970 444138 631977
rect 444354 632011 444562 632064
rect 444354 631977 444366 632011
rect 444550 631977 444562 632011
rect 444354 631970 444562 631977
rect 444914 632318 445122 632324
rect 444914 632064 445040 632318
rect 445092 632064 445122 632318
rect 444914 632017 445122 632064
rect 445474 632318 445682 632324
rect 445474 632064 445600 632318
rect 445652 632064 445682 632318
rect 445474 632017 445682 632064
rect 444914 632011 445134 632017
rect 444914 631977 444938 632011
rect 445122 631977 445134 632011
rect 444914 631971 445134 631977
rect 445474 632011 445706 632017
rect 445474 631977 445510 632011
rect 445694 631977 445706 632011
rect 445474 631971 445706 631977
rect 445936 632012 445970 632542
rect 446396 632478 446430 632542
rect 446370 632468 446442 632478
rect 446370 632364 446380 632468
rect 446432 632364 446442 632468
rect 446370 632354 446442 632364
rect 446508 632324 446542 632542
rect 446968 632478 447002 632542
rect 446942 632468 447014 632478
rect 446942 632364 446952 632468
rect 447004 632364 447014 632468
rect 446942 632354 447014 632364
rect 446494 632318 446558 632324
rect 446494 632064 446500 632318
rect 446552 632064 446558 632318
rect 446494 632058 446558 632064
rect 446072 632028 446292 632030
rect 446072 632017 446078 632028
rect 446070 632012 446078 632017
rect 445936 631972 446078 632012
rect 446286 632008 446292 632028
rect 444914 631970 445122 631971
rect 445474 631970 445682 631971
rect 443634 631918 443680 631970
rect 443634 629362 443640 631918
rect 443674 629362 443680 631918
rect 443634 629250 443680 629362
rect 444092 631918 444138 631970
rect 445936 631930 445970 631972
rect 446070 631971 446078 631972
rect 446072 631970 446078 631971
rect 446286 631972 446382 632008
rect 446286 631970 446292 631972
rect 446072 631960 446292 631970
rect 446508 631930 446542 632058
rect 446644 632024 446864 632030
rect 446644 632017 446650 632024
rect 446642 631971 446650 632017
rect 446644 631966 446650 631971
rect 446858 631966 446864 632024
rect 446644 631960 446864 631966
rect 447080 632012 447114 632542
rect 447540 632478 447574 632542
rect 447514 632468 447586 632478
rect 447514 632364 447524 632468
rect 447576 632364 447586 632468
rect 447514 632354 447586 632364
rect 447652 632324 447686 632542
rect 448112 632478 448146 632542
rect 448086 632468 448158 632478
rect 448086 632364 448096 632468
rect 448148 632364 448158 632468
rect 448086 632354 448158 632364
rect 447638 632318 447702 632324
rect 447638 632064 447644 632318
rect 447696 632064 447702 632318
rect 447638 632058 447702 632064
rect 447216 632028 447436 632034
rect 447216 632017 447222 632028
rect 447214 632012 447222 632017
rect 447080 631976 447222 632012
rect 447430 632012 447436 632028
rect 447080 631930 447114 631976
rect 447214 631971 447222 631976
rect 447216 631970 447222 631971
rect 447430 631976 447526 632012
rect 447430 631970 447436 631976
rect 447216 631964 447436 631970
rect 447652 631930 447686 632058
rect 447788 632028 448008 632034
rect 447788 632017 447794 632028
rect 447786 631971 447794 632017
rect 447788 631970 447794 631971
rect 448002 631970 448008 632028
rect 447788 631964 448008 631970
rect 448224 632012 448258 632542
rect 448684 632478 448718 632542
rect 448658 632468 448730 632478
rect 448658 632364 448668 632468
rect 448720 632364 448730 632468
rect 448658 632354 448730 632364
rect 448796 632324 448830 632542
rect 449256 632478 449290 632542
rect 449230 632468 449302 632478
rect 449230 632364 449240 632468
rect 449292 632364 449302 632468
rect 449230 632354 449302 632364
rect 448782 632318 448846 632324
rect 448782 632064 448788 632318
rect 448840 632064 448846 632318
rect 448782 632058 448846 632064
rect 449502 632318 449710 632324
rect 449502 632064 449588 632318
rect 449640 632064 449710 632318
rect 448360 632028 448580 632034
rect 448360 632017 448366 632028
rect 448358 632012 448366 632017
rect 448224 631976 448366 632012
rect 448574 632012 448580 632028
rect 448224 631930 448258 631976
rect 448358 631971 448366 631976
rect 448360 631970 448366 631971
rect 448574 631976 448670 632012
rect 448574 631970 448580 631976
rect 448360 631964 448580 631970
rect 448796 631930 448830 632058
rect 448932 632028 449152 632034
rect 448932 632017 448938 632028
rect 448930 631971 448938 632017
rect 448932 631970 448938 631971
rect 449146 631970 449152 632028
rect 449502 632011 449710 632064
rect 449502 631977 449514 632011
rect 449698 631977 449710 632011
rect 449502 631970 449710 631977
rect 450062 632318 450270 632324
rect 450062 632064 450148 632318
rect 450200 632064 450270 632318
rect 450062 632017 450270 632064
rect 450622 632318 450830 635726
rect 451884 634554 452016 637794
rect 452340 634694 452472 638378
rect 453858 638684 455858 639098
rect 453858 638396 453864 638684
rect 455852 638396 455858 638684
rect 453858 637190 455858 638396
rect 456558 638084 458558 638096
rect 456558 637796 456564 638084
rect 458552 637796 458558 638084
rect 456558 637190 458558 637796
rect 453898 637128 453938 637190
rect 454818 637128 454858 637190
rect 455738 637128 455778 637190
rect 452340 634614 452346 634694
rect 452466 634614 452472 634694
rect 452340 634608 452472 634614
rect 453442 637116 453488 637128
rect 451884 634474 451890 634554
rect 452000 634474 452016 634554
rect 451884 634468 452016 634474
rect 450622 632064 450708 632318
rect 450760 632064 450830 632318
rect 450622 632017 450830 632064
rect 452752 632318 453232 632324
rect 452752 632064 452758 632318
rect 453226 632064 453232 632318
rect 450062 632011 450282 632017
rect 450062 631977 450086 632011
rect 450270 631977 450282 632011
rect 450062 631971 450282 631977
rect 450622 632011 450854 632017
rect 450622 631977 450658 632011
rect 450842 631977 450854 632011
rect 450622 631971 450854 631977
rect 451070 632011 451574 632018
rect 451070 631977 451230 632011
rect 451414 631977 451574 632011
rect 450062 631970 450270 631971
rect 450622 631970 450830 631971
rect 451070 631970 451574 631977
rect 448932 631964 449152 631970
rect 444092 629362 444098 631918
rect 444132 629362 444138 631918
rect 444092 629250 444138 629362
rect 444206 631918 444252 631930
rect 444206 629362 444212 631918
rect 444246 629362 444252 631918
rect 444206 629350 444252 629362
rect 444664 631918 444710 631930
rect 444664 629362 444670 631918
rect 444704 629362 444710 631918
rect 444664 629350 444710 629362
rect 444778 631918 444824 631930
rect 444778 629362 444784 631918
rect 444818 629362 444824 631918
rect 444778 629350 444824 629362
rect 445236 631918 445282 631930
rect 445236 629362 445242 631918
rect 445276 631914 445282 631918
rect 445350 631918 445396 631930
rect 445276 629362 445284 631914
rect 445236 629350 445284 629362
rect 445350 629362 445356 631918
rect 445390 629362 445396 631918
rect 445350 629350 445396 629362
rect 445808 631918 445854 631930
rect 445808 629362 445814 631918
rect 445848 631914 445854 631918
rect 445922 631918 445970 631930
rect 445848 629362 445864 631914
rect 445808 629350 445864 629362
rect 445922 629362 445928 631918
rect 445962 631914 445970 631918
rect 446380 631918 446426 631930
rect 445962 629362 445968 631914
rect 445922 629350 445968 629362
rect 446380 629362 446386 631918
rect 446420 631914 446426 631918
rect 446494 631918 446542 631930
rect 446952 631918 446998 631930
rect 446420 629362 446428 631914
rect 446380 629350 446428 629362
rect 446494 629362 446500 631918
rect 446534 629362 446540 631918
rect 446494 629350 446540 629362
rect 446952 629362 446958 631918
rect 446992 631914 446998 631918
rect 447066 631918 447114 631930
rect 447524 631918 447570 631930
rect 446992 629362 447000 631914
rect 446952 629350 447000 629362
rect 447066 629362 447072 631918
rect 447106 629362 447112 631918
rect 447066 629350 447112 629362
rect 447524 629362 447530 631918
rect 447564 629362 447570 631918
rect 447524 629350 447570 629362
rect 447638 631918 447686 631930
rect 448096 631918 448142 631930
rect 447638 629362 447644 631918
rect 447678 629362 447684 631918
rect 447638 629350 447684 629362
rect 448096 629362 448102 631918
rect 448136 629362 448142 631918
rect 448096 629350 448142 629362
rect 448210 631918 448258 631930
rect 448668 631918 448714 631930
rect 448210 629362 448216 631918
rect 448250 629362 448256 631918
rect 448210 629350 448256 629362
rect 448668 629362 448674 631918
rect 448708 629362 448714 631918
rect 448668 629350 448714 629362
rect 448782 631918 448830 631930
rect 449240 631918 449286 631930
rect 448782 629362 448788 631918
rect 448822 629362 448828 631918
rect 448782 629350 448828 629362
rect 449240 629362 449246 631918
rect 449280 629362 449286 631918
rect 449240 629350 449286 629362
rect 449354 631918 449400 631930
rect 449354 629362 449360 631918
rect 449394 629362 449400 631918
rect 449354 629350 449400 629362
rect 449812 631918 449858 631930
rect 449812 629362 449818 631918
rect 449852 629362 449858 631918
rect 449812 629350 449858 629362
rect 449926 631918 449972 631930
rect 449926 629362 449932 631918
rect 449966 629362 449972 631918
rect 449926 629350 449972 629362
rect 450384 631918 450430 631930
rect 450384 629362 450390 631918
rect 450424 629362 450430 631918
rect 450384 629350 450430 629362
rect 450498 631918 450544 631930
rect 450498 629362 450504 631918
rect 450538 629362 450544 631918
rect 450498 629350 450544 629362
rect 450956 631918 451002 631930
rect 450956 629362 450962 631918
rect 450996 629362 451002 631918
rect 450956 629350 451002 629362
rect 451070 631918 451116 631970
rect 451070 629362 451076 631918
rect 451110 629362 451116 631918
rect 443620 629240 443692 629250
rect 443620 629136 443630 629240
rect 443682 629136 443692 629240
rect 443620 629126 443692 629136
rect 444078 629240 444150 629250
rect 444078 629136 444088 629240
rect 444140 629136 444150 629240
rect 444078 629126 444150 629136
rect 444208 629050 444250 629350
rect 444670 629250 444704 629350
rect 444654 629240 444726 629250
rect 444654 629136 444664 629240
rect 444716 629136 444726 629240
rect 444654 629126 444726 629136
rect 444780 629050 444822 629350
rect 445242 629250 445284 629350
rect 445226 629240 445298 629250
rect 445226 629136 445236 629240
rect 445288 629136 445298 629240
rect 445226 629126 445298 629136
rect 445352 629050 445394 629350
rect 445814 629250 445864 629350
rect 446386 629250 446428 629350
rect 446958 629250 447000 629350
rect 447530 629250 447564 629350
rect 448102 629250 448136 629350
rect 448674 629250 448708 629350
rect 449246 629250 449280 629350
rect 445798 629240 445870 629250
rect 445798 629136 445808 629240
rect 445860 629136 445870 629240
rect 445798 629126 445870 629136
rect 446370 629240 446442 629250
rect 446370 629136 446380 629240
rect 446432 629136 446442 629240
rect 446370 629126 446442 629136
rect 446942 629240 447014 629250
rect 446942 629136 446952 629240
rect 447004 629136 447014 629240
rect 446942 629126 447014 629136
rect 447514 629240 447586 629250
rect 447514 629136 447524 629240
rect 447576 629136 447586 629240
rect 447514 629126 447586 629136
rect 448086 629240 448158 629250
rect 448086 629136 448096 629240
rect 448148 629136 448158 629240
rect 448086 629126 448158 629136
rect 448658 629240 448730 629250
rect 448658 629136 448668 629240
rect 448720 629136 448730 629240
rect 448658 629126 448730 629136
rect 449230 629240 449298 629250
rect 449230 629136 449240 629240
rect 449292 629136 449298 629240
rect 449230 629126 449298 629136
rect 449356 629050 449398 629350
rect 449818 629250 449852 629350
rect 449802 629240 449870 629250
rect 449802 629136 449812 629240
rect 449864 629136 449870 629240
rect 449802 629126 449870 629136
rect 449928 629050 449970 629350
rect 450390 629250 450424 629350
rect 450374 629240 450442 629250
rect 450374 629136 450384 629240
rect 450436 629136 450442 629240
rect 450374 629126 450442 629136
rect 450500 629050 450542 629350
rect 450962 629250 450996 629350
rect 451070 629250 451116 629362
rect 451528 631918 451574 631970
rect 451528 629362 451534 631918
rect 451568 629362 451574 631918
rect 451528 629250 451574 629362
rect 452110 631830 452242 631842
rect 452110 629488 452126 631830
rect 452226 629488 452242 631830
rect 450946 629240 451014 629250
rect 450946 629136 450956 629240
rect 451008 629136 451014 629240
rect 450946 629126 451014 629136
rect 451056 629240 451128 629250
rect 451056 629136 451066 629240
rect 451118 629136 451128 629240
rect 451056 629126 451128 629136
rect 451514 629240 451586 629250
rect 451514 629136 451524 629240
rect 451576 629136 451586 629240
rect 451514 629126 451586 629136
rect 452110 629240 452242 629488
rect 452110 629136 452136 629240
rect 452188 629136 452242 629240
rect 452110 629126 452242 629136
rect 452752 629224 453232 632064
rect 452752 629076 452758 629224
rect 453226 629076 453232 629224
rect 452752 629070 453232 629076
rect 453442 629400 453448 637116
rect 453482 629400 453488 637116
rect 453898 637116 453946 637128
rect 453898 637090 453906 637116
rect 453442 629348 453488 629400
rect 453900 629400 453906 637090
rect 453940 629400 453946 637116
rect 453900 629384 453946 629400
rect 454358 637116 454404 637128
rect 454358 629400 454364 637116
rect 454398 629400 454404 637116
rect 454358 629388 454404 629400
rect 454816 637116 454862 637128
rect 454816 629400 454822 637116
rect 454856 629400 454862 637116
rect 454816 629388 454862 629400
rect 455274 637116 455320 637128
rect 455274 629400 455280 637116
rect 455314 629400 455320 637116
rect 455274 629388 455320 629400
rect 455732 637116 455778 637128
rect 455732 629400 455738 637116
rect 455772 629400 455778 637116
rect 455732 629388 455778 629400
rect 456190 637116 456236 637128
rect 456190 629400 456196 637116
rect 456230 629410 456236 637116
rect 456638 637116 456698 637190
rect 456638 637110 456654 637116
rect 456230 629400 456238 629410
rect 456190 629388 456238 629400
rect 456648 629400 456654 637110
rect 456688 637110 456698 637116
rect 457106 637116 457152 637128
rect 456688 629400 456694 637110
rect 457106 629410 457112 637116
rect 456648 629388 456694 629400
rect 457098 629400 457112 629410
rect 457146 629400 457152 637116
rect 457558 637116 457618 637190
rect 457558 637090 457570 637116
rect 457098 629388 457152 629400
rect 457564 629400 457570 637090
rect 457604 637090 457618 637116
rect 458022 637116 458068 637128
rect 457604 629400 457610 637090
rect 458022 629410 458028 637116
rect 457564 629388 457610 629400
rect 458018 629400 458028 629410
rect 458062 629400 458068 637116
rect 458478 637116 458538 637190
rect 459358 637188 464058 639982
rect 471526 640328 472474 640334
rect 471526 639810 471534 640328
rect 472468 639810 472474 640328
rect 467558 639548 469558 639590
rect 467558 639098 467564 639548
rect 469552 639098 469558 639548
rect 467558 638684 469558 639098
rect 467558 638396 467564 638684
rect 469552 638396 469558 638684
rect 464858 638084 466858 638096
rect 464858 637796 464864 638084
rect 466852 637796 466858 638084
rect 464858 637190 466858 637796
rect 467558 637190 469558 638396
rect 458478 637090 458486 637116
rect 458018 629388 458068 629400
rect 458480 629400 458486 637090
rect 458520 637090 458538 637116
rect 459398 637128 459438 637188
rect 460318 637128 460358 637188
rect 461238 637128 461278 637188
rect 462158 637128 462198 637188
rect 459398 637116 459446 637128
rect 459398 637110 459406 637116
rect 458520 629400 458526 637090
rect 458480 629388 458526 629400
rect 459400 629400 459406 637110
rect 459440 629400 459446 637116
rect 459400 629388 459446 629400
rect 459858 637116 459904 637128
rect 459858 629400 459864 637116
rect 459898 629400 459904 637116
rect 459858 629388 459904 629400
rect 460316 637116 460362 637128
rect 460316 629400 460322 637116
rect 460356 629400 460362 637116
rect 460316 629388 460362 629400
rect 460774 637116 460820 637128
rect 460774 629400 460780 637116
rect 460814 629400 460820 637116
rect 460774 629388 460820 629400
rect 461232 637116 461278 637128
rect 461232 629400 461238 637116
rect 461272 629400 461278 637116
rect 461232 629388 461278 629400
rect 461690 637116 461736 637128
rect 461690 629400 461696 637116
rect 461730 629410 461736 637116
rect 462148 637116 462198 637128
rect 461730 629400 461738 629410
rect 461690 629388 461738 629400
rect 462148 629400 462154 637116
rect 462188 637090 462198 637116
rect 462606 637116 462652 637128
rect 462188 629400 462194 637090
rect 462606 629410 462612 637116
rect 462148 629388 462194 629400
rect 462598 629400 462612 629410
rect 462646 629400 462652 637116
rect 463058 637116 463118 637188
rect 463058 637090 463070 637116
rect 462598 629388 462652 629400
rect 463064 629400 463070 637090
rect 463104 637090 463118 637116
rect 463522 637116 463568 637128
rect 463104 629400 463110 637090
rect 463522 629410 463528 637116
rect 463064 629388 463110 629400
rect 463518 629400 463528 629410
rect 463562 629400 463568 637116
rect 463978 637116 464038 637188
rect 463978 637090 463986 637116
rect 463518 629388 463568 629400
rect 463980 629400 463986 637090
rect 464020 637090 464038 637116
rect 464898 637128 464938 637190
rect 465818 637128 465858 637190
rect 466738 637128 466778 637190
rect 464898 637116 464946 637128
rect 464898 637090 464906 637116
rect 464020 629400 464026 637090
rect 463980 629388 464026 629400
rect 464900 629400 464906 637090
rect 464940 629400 464946 637116
rect 464900 629388 464946 629400
rect 465358 637116 465404 637128
rect 465358 629400 465364 637116
rect 465398 629400 465404 637116
rect 465358 629388 465404 629400
rect 465816 637116 465862 637128
rect 465816 629400 465822 637116
rect 465856 629400 465862 637116
rect 465816 629388 465862 629400
rect 466274 637116 466320 637128
rect 466274 629400 466280 637116
rect 466314 629400 466320 637116
rect 466274 629388 466320 629400
rect 466732 637116 466778 637128
rect 466732 629400 466738 637116
rect 466772 629400 466778 637116
rect 466732 629388 466778 629400
rect 467190 637116 467236 637128
rect 467190 629400 467196 637116
rect 467230 629410 467236 637116
rect 467638 637116 467698 637190
rect 467638 637090 467654 637116
rect 467230 629400 467238 629410
rect 467190 629388 467238 629400
rect 467648 629400 467654 637090
rect 467688 637090 467698 637116
rect 468106 637116 468152 637128
rect 467688 629400 467694 637090
rect 468106 629410 468112 637116
rect 467648 629388 467694 629400
rect 468098 629400 468112 629410
rect 468146 629400 468152 637116
rect 468558 637116 468618 637190
rect 469478 637128 469518 637190
rect 468558 637110 468570 637116
rect 468098 629388 468152 629400
rect 468564 629400 468570 637110
rect 468604 637110 468618 637116
rect 469022 637116 469068 637128
rect 468604 629400 468610 637110
rect 469022 629410 469028 637116
rect 468564 629388 468610 629400
rect 469018 629400 469028 629410
rect 469062 629400 469068 637116
rect 469478 637116 469526 637128
rect 469478 637110 469486 637116
rect 469018 629388 469068 629400
rect 469480 629400 469486 637110
rect 469520 629400 469526 637116
rect 453442 629347 453590 629348
rect 453782 629347 453900 629348
rect 454058 629347 454238 629350
rect 453442 629341 453900 629347
rect 453442 629307 453602 629341
rect 453786 629307 453900 629341
rect 443318 628932 443324 629046
rect 443518 628932 443524 629046
rect 443318 628926 443524 628932
rect 444194 629040 444266 629050
rect 444194 628936 444204 629040
rect 444256 628936 444266 629040
rect 444194 628926 444266 628936
rect 444766 629040 444838 629050
rect 444766 628936 444776 629040
rect 444828 628936 444838 629040
rect 444766 628926 444838 628936
rect 445338 629040 445410 629050
rect 445338 628936 445348 629040
rect 445400 628936 445410 629040
rect 449342 629040 449414 629050
rect 445338 628926 445410 628936
rect 446568 628984 449022 629000
rect 446568 628884 446580 628984
rect 448922 628884 449022 628984
rect 449342 628936 449352 629040
rect 449404 628936 449414 629040
rect 449342 628926 449414 628936
rect 449914 629040 449986 629050
rect 449914 628936 449924 629040
rect 449976 628936 449986 629040
rect 449914 628926 449986 628936
rect 450486 629040 450558 629050
rect 450486 628936 450496 629040
rect 450548 628936 450558 629040
rect 453442 628990 453900 629307
rect 454048 629341 454256 629347
rect 454048 629307 454060 629341
rect 454244 629307 454256 629341
rect 454048 629301 454256 629307
rect 454058 629210 454238 629301
rect 454058 629090 454078 629210
rect 454218 629090 454238 629210
rect 454058 629070 454238 629090
rect 454358 629030 454398 629388
rect 454518 629347 454698 629350
rect 454978 629347 455158 629350
rect 454506 629341 454714 629347
rect 454506 629307 454518 629341
rect 454702 629307 454714 629341
rect 454506 629301 454714 629307
rect 454964 629341 455172 629347
rect 454964 629307 454976 629341
rect 455160 629307 455172 629341
rect 454964 629301 455172 629307
rect 454518 629210 454698 629301
rect 454518 629090 454538 629210
rect 454678 629090 454698 629210
rect 454518 629070 454698 629090
rect 454978 629210 455158 629301
rect 454978 629090 454998 629210
rect 455138 629090 455158 629210
rect 454978 629070 455158 629090
rect 455278 629030 455318 629388
rect 455438 629347 455618 629350
rect 455898 629347 456078 629350
rect 455422 629341 455630 629347
rect 455422 629307 455434 629341
rect 455618 629307 455630 629341
rect 455422 629301 455630 629307
rect 455880 629341 456088 629347
rect 455880 629307 455892 629341
rect 456076 629307 456088 629341
rect 455880 629301 456088 629307
rect 455438 629210 455618 629301
rect 455438 629090 455458 629210
rect 455598 629090 455618 629210
rect 455438 629070 455618 629090
rect 455898 629210 456078 629301
rect 455898 629090 455918 629210
rect 456058 629090 456078 629210
rect 455898 629070 456078 629090
rect 456198 629030 456238 629388
rect 456358 629347 456538 629350
rect 456818 629347 456998 629350
rect 456338 629341 456546 629347
rect 456338 629307 456350 629341
rect 456534 629307 456546 629341
rect 456338 629301 456546 629307
rect 456796 629341 457004 629347
rect 456796 629307 456808 629341
rect 456992 629307 457004 629341
rect 456796 629301 457004 629307
rect 456358 629210 456538 629301
rect 456358 629090 456378 629210
rect 456518 629090 456538 629210
rect 456358 629070 456538 629090
rect 456818 629210 456998 629301
rect 456818 629090 456838 629210
rect 456978 629090 456998 629210
rect 456818 629070 456998 629090
rect 457098 629030 457138 629388
rect 457278 629347 457458 629350
rect 457738 629347 457918 629350
rect 457254 629341 457462 629347
rect 457254 629307 457266 629341
rect 457450 629307 457462 629341
rect 457254 629301 457462 629307
rect 457712 629341 457920 629347
rect 457712 629307 457724 629341
rect 457908 629307 457920 629341
rect 457712 629301 457920 629307
rect 457278 629210 457458 629301
rect 457278 629090 457298 629210
rect 457438 629090 457458 629210
rect 457278 629070 457458 629090
rect 457738 629210 457918 629301
rect 457738 629090 457758 629210
rect 457898 629090 457918 629210
rect 457738 629070 457918 629090
rect 458018 629030 458058 629388
rect 458198 629347 458378 629350
rect 459558 629347 459738 629350
rect 458170 629341 458378 629347
rect 458170 629307 458182 629341
rect 458366 629307 458378 629341
rect 458170 629301 458378 629307
rect 459548 629341 459756 629347
rect 459548 629307 459560 629341
rect 459744 629307 459756 629341
rect 459548 629301 459756 629307
rect 458198 629210 458378 629301
rect 458198 629090 458218 629210
rect 458358 629090 458378 629210
rect 458198 629070 458378 629090
rect 459558 629210 459738 629301
rect 459558 629090 459578 629210
rect 459718 629090 459738 629210
rect 459558 629070 459738 629090
rect 459858 629030 459898 629388
rect 460018 629347 460198 629350
rect 460478 629347 460658 629350
rect 460006 629341 460214 629347
rect 460006 629307 460018 629341
rect 460202 629307 460214 629341
rect 460006 629301 460214 629307
rect 460464 629341 460672 629347
rect 460464 629307 460476 629341
rect 460660 629307 460672 629341
rect 460464 629301 460672 629307
rect 460018 629210 460198 629301
rect 460018 629090 460038 629210
rect 460178 629090 460198 629210
rect 460018 629070 460198 629090
rect 460478 629210 460658 629301
rect 460478 629090 460498 629210
rect 460638 629090 460658 629210
rect 460478 629070 460658 629090
rect 460778 629030 460818 629388
rect 460938 629347 461118 629350
rect 461398 629347 461578 629350
rect 460922 629341 461130 629347
rect 460922 629307 460934 629341
rect 461118 629307 461130 629341
rect 460922 629301 461130 629307
rect 461380 629341 461588 629347
rect 461380 629307 461392 629341
rect 461576 629307 461588 629341
rect 461380 629301 461588 629307
rect 460938 629210 461118 629301
rect 460938 629090 460958 629210
rect 461098 629090 461118 629210
rect 460938 629070 461118 629090
rect 461398 629210 461578 629301
rect 461398 629090 461418 629210
rect 461558 629090 461578 629210
rect 461398 629070 461578 629090
rect 461698 629030 461738 629388
rect 461858 629347 462038 629350
rect 462318 629347 462498 629350
rect 461838 629341 462046 629347
rect 461838 629307 461850 629341
rect 462034 629307 462046 629341
rect 461838 629301 462046 629307
rect 462296 629341 462504 629347
rect 462296 629307 462308 629341
rect 462492 629307 462504 629341
rect 462296 629301 462504 629307
rect 461858 629210 462038 629301
rect 461858 629090 461878 629210
rect 462018 629090 462038 629210
rect 461858 629070 462038 629090
rect 462318 629210 462498 629301
rect 462318 629090 462338 629210
rect 462478 629090 462498 629210
rect 462318 629070 462498 629090
rect 462598 629030 462638 629388
rect 462778 629347 462958 629350
rect 463238 629347 463418 629350
rect 462754 629341 462962 629347
rect 462754 629307 462766 629341
rect 462950 629307 462962 629341
rect 462754 629301 462962 629307
rect 463212 629341 463420 629347
rect 463212 629307 463224 629341
rect 463408 629307 463420 629341
rect 463212 629301 463420 629307
rect 462778 629210 462958 629301
rect 462778 629090 462798 629210
rect 462938 629090 462958 629210
rect 462778 629070 462958 629090
rect 463238 629210 463418 629301
rect 463238 629090 463258 629210
rect 463398 629090 463418 629210
rect 463238 629070 463418 629090
rect 463518 629030 463558 629388
rect 463698 629347 463878 629350
rect 465058 629347 465238 629350
rect 463670 629341 463878 629347
rect 463670 629307 463682 629341
rect 463866 629307 463878 629341
rect 463670 629301 463878 629307
rect 465048 629341 465256 629347
rect 465048 629307 465060 629341
rect 465244 629307 465256 629341
rect 465048 629301 465256 629307
rect 463698 629210 463878 629301
rect 463698 629090 463718 629210
rect 463858 629090 463878 629210
rect 463698 629070 463878 629090
rect 465058 629210 465238 629301
rect 465058 629090 465078 629210
rect 465218 629090 465238 629210
rect 465058 629070 465238 629090
rect 465358 629030 465398 629388
rect 465518 629347 465698 629350
rect 465978 629347 466158 629350
rect 465506 629341 465714 629347
rect 465506 629307 465518 629341
rect 465702 629307 465714 629341
rect 465506 629301 465714 629307
rect 465964 629341 466172 629347
rect 465964 629307 465976 629341
rect 466160 629307 466172 629341
rect 465964 629301 466172 629307
rect 465518 629210 465698 629301
rect 465518 629090 465538 629210
rect 465678 629090 465698 629210
rect 465518 629070 465698 629090
rect 465978 629210 466158 629301
rect 465978 629090 465998 629210
rect 466138 629090 466158 629210
rect 465978 629070 466158 629090
rect 466278 629030 466318 629388
rect 466438 629347 466618 629350
rect 466898 629347 467078 629350
rect 466422 629341 466630 629347
rect 466422 629307 466434 629341
rect 466618 629307 466630 629341
rect 466422 629301 466630 629307
rect 466880 629341 467088 629347
rect 466880 629307 466892 629341
rect 467076 629307 467088 629341
rect 466880 629301 467088 629307
rect 466438 629210 466618 629301
rect 466438 629090 466458 629210
rect 466598 629090 466618 629210
rect 466438 629070 466618 629090
rect 466898 629210 467078 629301
rect 466898 629090 466918 629210
rect 467058 629090 467078 629210
rect 466898 629070 467078 629090
rect 467198 629030 467238 629388
rect 467358 629347 467538 629350
rect 467818 629347 467998 629350
rect 467338 629341 467546 629347
rect 467338 629307 467350 629341
rect 467534 629307 467546 629341
rect 467338 629301 467546 629307
rect 467796 629341 468004 629347
rect 467796 629307 467808 629341
rect 467992 629307 468004 629341
rect 467796 629301 468004 629307
rect 467358 629210 467538 629301
rect 467358 629090 467378 629210
rect 467518 629090 467538 629210
rect 467358 629070 467538 629090
rect 467818 629210 467998 629301
rect 467818 629090 467838 629210
rect 467978 629090 467998 629210
rect 467818 629070 467998 629090
rect 468098 629030 468138 629388
rect 468278 629347 468458 629350
rect 468738 629347 468918 629350
rect 468254 629341 468462 629347
rect 468254 629307 468266 629341
rect 468450 629307 468462 629341
rect 468254 629301 468462 629307
rect 468712 629341 468920 629347
rect 468712 629307 468724 629341
rect 468908 629307 468920 629341
rect 468712 629301 468920 629307
rect 468278 629210 468458 629301
rect 468278 629090 468298 629210
rect 468438 629090 468458 629210
rect 468278 629070 468458 629090
rect 468738 629210 468918 629301
rect 468738 629090 468758 629210
rect 468898 629090 468918 629210
rect 468738 629070 468918 629090
rect 469018 629030 469058 629388
rect 469480 629384 469526 629400
rect 469938 637116 469984 637128
rect 469938 629400 469944 637116
rect 469978 629400 469984 637116
rect 471526 630850 472474 639810
rect 472870 639548 473574 642186
rect 472870 639098 472876 639548
rect 473568 639098 473574 639548
rect 472870 635760 473574 639098
rect 473688 642878 474392 642884
rect 473688 642186 473694 642878
rect 474386 642186 474392 642878
rect 474588 642867 475150 642873
rect 474588 642470 474600 642867
rect 475138 642470 475150 642867
rect 474588 642464 475150 642470
rect 473688 638084 474392 642186
rect 475667 638987 480819 639597
rect 473688 637796 473696 638084
rect 474386 637796 474392 638084
rect 473688 637790 474392 637796
rect 475057 636999 480819 638987
rect 475667 636411 480819 636999
rect 472870 635068 472876 635760
rect 473568 635068 473574 635760
rect 472870 635060 473574 635068
rect 471526 629914 471532 630850
rect 472468 629914 472474 630850
rect 475057 634445 476955 636411
rect 478921 634445 480819 636411
rect 475057 630550 480819 634445
rect 475057 630498 476352 630550
rect 476404 630498 476456 630550
rect 476508 630498 476560 630550
rect 476612 630498 476664 630550
rect 476716 630498 476768 630550
rect 476820 630498 476872 630550
rect 476924 630498 480819 630550
rect 475057 630446 480819 630498
rect 475057 630394 476352 630446
rect 476404 630394 476456 630446
rect 476508 630394 476560 630446
rect 476612 630394 476664 630446
rect 476716 630394 476768 630446
rect 476820 630394 476872 630446
rect 476924 630394 480819 630446
rect 475057 630342 480819 630394
rect 475057 630290 476352 630342
rect 476404 630290 476456 630342
rect 476508 630290 476560 630342
rect 476612 630290 476664 630342
rect 476716 630290 476768 630342
rect 476820 630290 476872 630342
rect 476924 630290 480819 630342
rect 475057 630238 480819 630290
rect 475057 630186 476352 630238
rect 476404 630186 476456 630238
rect 476508 630186 476560 630238
rect 476612 630186 476664 630238
rect 476716 630186 476768 630238
rect 476820 630186 476872 630238
rect 476924 630186 480819 630238
rect 475057 630134 480819 630186
rect 482144 636778 483202 636788
rect 482144 636678 482174 636778
rect 482274 636678 482398 636778
rect 482498 636678 482622 636778
rect 482722 636678 482846 636778
rect 482946 636678 483070 636778
rect 483170 636678 483202 636778
rect 482144 636554 483202 636678
rect 482144 636454 482174 636554
rect 482274 636454 482398 636554
rect 482498 636454 482622 636554
rect 482722 636454 482846 636554
rect 482946 636454 483070 636554
rect 483170 636454 483202 636554
rect 482144 636330 483202 636454
rect 482144 636230 482174 636330
rect 482274 636230 482398 636330
rect 482498 636230 482622 636330
rect 482722 636230 482846 636330
rect 482946 636230 483070 636330
rect 483170 636230 483202 636330
rect 482144 636106 483202 636230
rect 482144 636006 482174 636106
rect 482274 636006 482398 636106
rect 482498 636006 482622 636106
rect 482722 636006 482846 636106
rect 482946 636006 483070 636106
rect 483170 636006 483202 636106
rect 482144 635882 483202 636006
rect 482144 635782 482174 635882
rect 482274 635782 482398 635882
rect 482498 635782 482622 635882
rect 482722 635782 482846 635882
rect 482946 635782 483070 635882
rect 483170 635782 483202 635882
rect 482144 635658 483202 635782
rect 482144 635558 482174 635658
rect 482274 635558 482398 635658
rect 482498 635558 482622 635658
rect 482722 635558 482846 635658
rect 482946 635558 483070 635658
rect 483170 635558 483202 635658
rect 482144 635434 483202 635558
rect 482144 635334 482174 635434
rect 482274 635334 482398 635434
rect 482498 635334 482622 635434
rect 482722 635334 482846 635434
rect 482946 635334 483070 635434
rect 483170 635334 483202 635434
rect 482144 635210 483202 635334
rect 482144 635110 482174 635210
rect 482274 635110 482398 635210
rect 482498 635110 482622 635210
rect 482722 635110 482846 635210
rect 482946 635110 483070 635210
rect 483170 635110 483202 635210
rect 482144 634986 483202 635110
rect 482144 634886 482174 634986
rect 482274 634886 482398 634986
rect 482498 634886 482622 634986
rect 482722 634886 482846 634986
rect 482946 634886 483070 634986
rect 483170 634886 483202 634986
rect 482144 634762 483202 634886
rect 482144 634662 482174 634762
rect 482274 634662 482398 634762
rect 482498 634662 482622 634762
rect 482722 634662 482846 634762
rect 482946 634662 483070 634762
rect 483170 634662 483202 634762
rect 482144 634538 483202 634662
rect 482144 634438 482174 634538
rect 482274 634438 482398 634538
rect 482498 634438 482622 634538
rect 482722 634438 482846 634538
rect 482946 634438 483070 634538
rect 483170 634438 483202 634538
rect 482144 634314 483202 634438
rect 482144 634214 482174 634314
rect 482274 634214 482398 634314
rect 482498 634214 482622 634314
rect 482722 634214 482846 634314
rect 482946 634214 483070 634314
rect 483170 634214 483202 634314
rect 482144 634090 483202 634214
rect 482144 633990 482174 634090
rect 482274 633990 482398 634090
rect 482498 633990 482622 634090
rect 482722 633990 482846 634090
rect 482946 633990 483070 634090
rect 483170 633990 483202 634090
rect 482144 633866 483202 633990
rect 482144 633766 482174 633866
rect 482274 633766 482398 633866
rect 482498 633766 482622 633866
rect 482722 633766 482846 633866
rect 482946 633766 483070 633866
rect 483170 633766 483202 633866
rect 482144 633642 483202 633766
rect 482144 633542 482174 633642
rect 482274 633542 482398 633642
rect 482498 633542 482622 633642
rect 482722 633542 482846 633642
rect 482946 633542 483070 633642
rect 483170 633542 483202 633642
rect 482144 633418 483202 633542
rect 482144 633318 482174 633418
rect 482274 633318 482398 633418
rect 482498 633318 482622 633418
rect 482722 633318 482846 633418
rect 482946 633318 483070 633418
rect 483170 633318 483202 633418
rect 482144 633194 483202 633318
rect 482144 633094 482174 633194
rect 482274 633094 482398 633194
rect 482498 633094 482622 633194
rect 482722 633094 482846 633194
rect 482946 633094 483070 633194
rect 483170 633094 483202 633194
rect 482144 632970 483202 633094
rect 482144 632870 482174 632970
rect 482274 632870 482398 632970
rect 482498 632870 482622 632970
rect 482722 632870 482846 632970
rect 482946 632870 483070 632970
rect 483170 632870 483202 632970
rect 482144 632746 483202 632870
rect 482144 632646 482174 632746
rect 482274 632646 482398 632746
rect 482498 632646 482622 632746
rect 482722 632646 482846 632746
rect 482946 632646 483070 632746
rect 483170 632646 483202 632746
rect 482144 632522 483202 632646
rect 482144 632422 482174 632522
rect 482274 632422 482398 632522
rect 482498 632422 482622 632522
rect 482722 632422 482846 632522
rect 482946 632422 483070 632522
rect 483170 632422 483202 632522
rect 482144 632298 483202 632422
rect 482144 632198 482174 632298
rect 482274 632198 482398 632298
rect 482498 632198 482622 632298
rect 482722 632198 482846 632298
rect 482946 632198 483070 632298
rect 483170 632198 483202 632298
rect 482144 632074 483202 632198
rect 482144 631974 482174 632074
rect 482274 631974 482398 632074
rect 482498 631974 482622 632074
rect 482722 631974 482846 632074
rect 482946 631974 483070 632074
rect 483170 631974 483202 632074
rect 482144 631850 483202 631974
rect 482144 631750 482174 631850
rect 482274 631750 482398 631850
rect 482498 631750 482622 631850
rect 482722 631750 482846 631850
rect 482946 631750 483070 631850
rect 483170 631750 483202 631850
rect 482144 631626 483202 631750
rect 482144 631526 482174 631626
rect 482274 631526 482398 631626
rect 482498 631526 482622 631626
rect 482722 631526 482846 631626
rect 482946 631526 483070 631626
rect 483170 631526 483202 631626
rect 482144 631402 483202 631526
rect 482144 631302 482174 631402
rect 482274 631302 482398 631402
rect 482498 631302 482622 631402
rect 482722 631302 482846 631402
rect 482946 631302 483070 631402
rect 483170 631302 483202 631402
rect 482144 631178 483202 631302
rect 482144 631078 482174 631178
rect 482274 631078 482398 631178
rect 482498 631078 482622 631178
rect 482722 631078 482846 631178
rect 482946 631078 483070 631178
rect 483170 631078 483202 631178
rect 482144 630954 483202 631078
rect 482144 630854 482174 630954
rect 482274 630854 482398 630954
rect 482498 630854 482622 630954
rect 482722 630854 482846 630954
rect 482946 630854 483070 630954
rect 483170 630854 483202 630954
rect 482144 630730 483202 630854
rect 482144 630630 482174 630730
rect 482274 630630 482398 630730
rect 482498 630630 482622 630730
rect 482722 630630 482846 630730
rect 482946 630630 483070 630730
rect 483170 630630 483202 630730
rect 482144 630506 483202 630630
rect 482144 630406 482174 630506
rect 482274 630406 482398 630506
rect 482498 630406 482622 630506
rect 482722 630406 482846 630506
rect 482946 630406 483070 630506
rect 483170 630406 483202 630506
rect 482144 630282 483202 630406
rect 482144 630182 482174 630282
rect 482274 630182 482398 630282
rect 482498 630182 482622 630282
rect 482722 630182 482846 630282
rect 482946 630182 483070 630282
rect 483170 630182 483202 630282
rect 482144 630162 483202 630182
rect 475057 630082 476352 630134
rect 476404 630082 476456 630134
rect 476508 630082 476560 630134
rect 476612 630082 476664 630134
rect 476716 630082 476768 630134
rect 476820 630082 476872 630134
rect 476924 630082 480819 630134
rect 475057 630030 480819 630082
rect 475057 629978 476352 630030
rect 476404 629978 476456 630030
rect 476508 629978 476560 630030
rect 476612 629978 476664 630030
rect 476716 629978 476768 630030
rect 476820 629978 476872 630030
rect 476924 629978 480819 630030
rect 475057 629971 480819 629978
rect 471526 629908 472474 629914
rect 469198 629347 469378 629350
rect 469938 629348 469984 629400
rect 469170 629341 469378 629347
rect 469170 629307 469182 629341
rect 469366 629307 469378 629341
rect 469170 629301 469378 629307
rect 469198 629210 469378 629301
rect 469198 629090 469218 629210
rect 469358 629090 469378 629210
rect 469198 629070 469378 629090
rect 469526 629341 469984 629348
rect 469526 629307 469640 629341
rect 469824 629307 469984 629341
rect 450486 628926 450558 628936
rect 446568 628868 449022 628884
rect 452748 628890 453900 628990
rect 454318 629010 454438 629030
rect 454318 628930 454338 629010
rect 454418 628930 454438 629010
rect 454318 628910 454438 628930
rect 455238 629010 455358 629030
rect 455238 628930 455258 629010
rect 455338 628930 455358 629010
rect 455238 628910 455358 628930
rect 456158 629010 456278 629030
rect 456158 628930 456178 629010
rect 456258 628930 456278 629010
rect 456158 628910 456278 628930
rect 457078 629010 457198 629030
rect 457078 628930 457098 629010
rect 457178 628930 457198 629010
rect 457078 628910 457198 628930
rect 457998 629010 458118 629030
rect 457998 628930 458018 629010
rect 458098 628930 458118 629010
rect 459818 629010 459938 629030
rect 457998 628910 458118 628930
rect 452748 628790 452848 628890
rect 453248 628790 453900 628890
rect 452748 628690 453900 628790
rect 458658 628890 459258 628990
rect 459818 628930 459838 629010
rect 459918 628930 459938 629010
rect 459818 628910 459938 628930
rect 460738 629010 460858 629030
rect 460738 628930 460758 629010
rect 460838 628930 460858 629010
rect 460738 628910 460858 628930
rect 461658 629010 461778 629030
rect 461658 628930 461678 629010
rect 461758 628930 461778 629010
rect 461658 628910 461778 628930
rect 462578 629010 462698 629030
rect 462578 628930 462598 629010
rect 462678 628930 462698 629010
rect 462578 628910 462698 628930
rect 463498 629010 463618 629030
rect 463498 628930 463518 629010
rect 463598 628930 463618 629010
rect 465318 629010 465438 629030
rect 463498 628910 463618 628930
rect 458658 628790 458758 628890
rect 459158 628790 459258 628890
rect 458658 628690 459258 628790
rect 464158 628890 464758 628990
rect 465318 628930 465338 629010
rect 465418 628930 465438 629010
rect 465318 628910 465438 628930
rect 466238 629010 466358 629030
rect 466238 628930 466258 629010
rect 466338 628930 466358 629010
rect 466238 628910 466358 628930
rect 467158 629010 467278 629030
rect 467158 628930 467178 629010
rect 467258 628930 467278 629010
rect 467158 628910 467278 628930
rect 468078 629010 468198 629030
rect 468078 628930 468098 629010
rect 468178 628930 468198 629010
rect 468078 628910 468198 628930
rect 468998 629010 469118 629030
rect 468998 628930 469018 629010
rect 469098 628930 469118 629010
rect 468998 628910 469118 628930
rect 469526 628988 469984 629307
rect 464158 628790 464258 628890
rect 464658 628790 464758 628890
rect 464158 628690 464758 628790
rect 469526 628888 470714 628988
rect 469526 628788 470214 628888
rect 470614 628788 470714 628888
rect 469526 628688 470714 628788
rect 438880 627656 445540 627686
rect 438880 627556 438920 627656
rect 439020 627556 439144 627656
rect 439244 627556 439368 627656
rect 439468 627556 439592 627656
rect 439692 627556 439816 627656
rect 439916 627556 440040 627656
rect 440140 627556 440264 627656
rect 440364 627556 440488 627656
rect 440588 627556 440712 627656
rect 440812 627556 440936 627656
rect 441036 627556 441160 627656
rect 441260 627556 441384 627656
rect 441484 627556 441608 627656
rect 441708 627556 441832 627656
rect 441932 627556 442056 627656
rect 442156 627556 442280 627656
rect 442380 627556 442504 627656
rect 442604 627556 442728 627656
rect 442828 627556 442952 627656
rect 443052 627556 443176 627656
rect 443276 627556 443400 627656
rect 443500 627556 443624 627656
rect 443724 627556 443848 627656
rect 443948 627556 444072 627656
rect 444172 627556 444296 627656
rect 444396 627556 444520 627656
rect 444620 627556 444744 627656
rect 444844 627556 444968 627656
rect 445068 627556 445192 627656
rect 445292 627556 445416 627656
rect 445516 627556 445540 627656
rect 438880 627432 445540 627556
rect 438880 627332 438920 627432
rect 439020 627332 439144 627432
rect 439244 627332 439368 627432
rect 439468 627332 439592 627432
rect 439692 627332 439816 627432
rect 439916 627332 440040 627432
rect 440140 627332 440264 627432
rect 440364 627332 440488 627432
rect 440588 627332 440712 627432
rect 440812 627332 440936 627432
rect 441036 627332 441160 627432
rect 441260 627332 441384 627432
rect 441484 627332 441608 627432
rect 441708 627332 441832 627432
rect 441932 627332 442056 627432
rect 442156 627332 442280 627432
rect 442380 627332 442504 627432
rect 442604 627332 442728 627432
rect 442828 627332 442952 627432
rect 443052 627332 443176 627432
rect 443276 627332 443400 627432
rect 443500 627332 443624 627432
rect 443724 627332 443848 627432
rect 443948 627332 444072 627432
rect 444172 627332 444296 627432
rect 444396 627332 444520 627432
rect 444620 627332 444744 627432
rect 444844 627332 444968 627432
rect 445068 627332 445192 627432
rect 445292 627332 445416 627432
rect 445516 627332 445540 627432
rect 438880 627208 445540 627332
rect 438880 627108 438920 627208
rect 439020 627108 439144 627208
rect 439244 627108 439368 627208
rect 439468 627108 439592 627208
rect 439692 627108 439816 627208
rect 439916 627108 440040 627208
rect 440140 627108 440264 627208
rect 440364 627108 440488 627208
rect 440588 627108 440712 627208
rect 440812 627108 440936 627208
rect 441036 627108 441160 627208
rect 441260 627108 441384 627208
rect 441484 627108 441608 627208
rect 441708 627108 441832 627208
rect 441932 627108 442056 627208
rect 442156 627108 442280 627208
rect 442380 627108 442504 627208
rect 442604 627108 442728 627208
rect 442828 627108 442952 627208
rect 443052 627108 443176 627208
rect 443276 627108 443400 627208
rect 443500 627108 443624 627208
rect 443724 627108 443848 627208
rect 443948 627108 444072 627208
rect 444172 627108 444296 627208
rect 444396 627108 444520 627208
rect 444620 627108 444744 627208
rect 444844 627108 444968 627208
rect 445068 627108 445192 627208
rect 445292 627108 445416 627208
rect 445516 627108 445540 627208
rect 438880 626984 445540 627108
rect 438880 626884 438920 626984
rect 439020 626884 439144 626984
rect 439244 626884 439368 626984
rect 439468 626884 439592 626984
rect 439692 626884 439816 626984
rect 439916 626884 440040 626984
rect 440140 626884 440264 626984
rect 440364 626884 440488 626984
rect 440588 626884 440712 626984
rect 440812 626884 440936 626984
rect 441036 626884 441160 626984
rect 441260 626884 441384 626984
rect 441484 626884 441608 626984
rect 441708 626884 441832 626984
rect 441932 626884 442056 626984
rect 442156 626884 442280 626984
rect 442380 626884 442504 626984
rect 442604 626884 442728 626984
rect 442828 626884 442952 626984
rect 443052 626884 443176 626984
rect 443276 626884 443400 626984
rect 443500 626884 443624 626984
rect 443724 626884 443848 626984
rect 443948 626884 444072 626984
rect 444172 626884 444296 626984
rect 444396 626884 444520 626984
rect 444620 626884 444744 626984
rect 444844 626884 444968 626984
rect 445068 626884 445192 626984
rect 445292 626884 445416 626984
rect 445516 626884 445540 626984
rect 438880 626760 445540 626884
rect 438880 626660 438920 626760
rect 439020 626660 439144 626760
rect 439244 626660 439368 626760
rect 439468 626660 439592 626760
rect 439692 626660 439816 626760
rect 439916 626660 440040 626760
rect 440140 626660 440264 626760
rect 440364 626660 440488 626760
rect 440588 626660 440712 626760
rect 440812 626660 440936 626760
rect 441036 626660 441160 626760
rect 441260 626660 441384 626760
rect 441484 626660 441608 626760
rect 441708 626660 441832 626760
rect 441932 626660 442056 626760
rect 442156 626660 442280 626760
rect 442380 626660 442504 626760
rect 442604 626660 442728 626760
rect 442828 626660 442952 626760
rect 443052 626660 443176 626760
rect 443276 626660 443400 626760
rect 443500 626660 443624 626760
rect 443724 626660 443848 626760
rect 443948 626660 444072 626760
rect 444172 626660 444296 626760
rect 444396 626660 444520 626760
rect 444620 626660 444744 626760
rect 444844 626660 444968 626760
rect 445068 626660 445192 626760
rect 445292 626660 445416 626760
rect 445516 626660 445540 626760
rect 438880 626626 445540 626660
rect 449350 627656 456010 627686
rect 449350 627556 449390 627656
rect 449490 627556 449614 627656
rect 449714 627556 449838 627656
rect 449938 627556 450062 627656
rect 450162 627556 450286 627656
rect 450386 627556 450510 627656
rect 450610 627556 450734 627656
rect 450834 627556 450958 627656
rect 451058 627556 451182 627656
rect 451282 627556 451406 627656
rect 451506 627556 451630 627656
rect 451730 627556 451854 627656
rect 451954 627556 452078 627656
rect 452178 627556 452302 627656
rect 452402 627556 452526 627656
rect 452626 627556 452750 627656
rect 452850 627556 452974 627656
rect 453074 627556 453198 627656
rect 453298 627556 453422 627656
rect 453522 627556 453646 627656
rect 453746 627556 453870 627656
rect 453970 627556 454094 627656
rect 454194 627556 454318 627656
rect 454418 627556 454542 627656
rect 454642 627556 454766 627656
rect 454866 627556 454990 627656
rect 455090 627556 455214 627656
rect 455314 627556 455438 627656
rect 455538 627556 455662 627656
rect 455762 627556 455886 627656
rect 455986 627556 456010 627656
rect 449350 627432 456010 627556
rect 449350 627332 449390 627432
rect 449490 627332 449614 627432
rect 449714 627332 449838 627432
rect 449938 627332 450062 627432
rect 450162 627332 450286 627432
rect 450386 627332 450510 627432
rect 450610 627332 450734 627432
rect 450834 627332 450958 627432
rect 451058 627332 451182 627432
rect 451282 627332 451406 627432
rect 451506 627332 451630 627432
rect 451730 627332 451854 627432
rect 451954 627332 452078 627432
rect 452178 627332 452302 627432
rect 452402 627332 452526 627432
rect 452626 627332 452750 627432
rect 452850 627332 452974 627432
rect 453074 627332 453198 627432
rect 453298 627332 453422 627432
rect 453522 627332 453646 627432
rect 453746 627332 453870 627432
rect 453970 627332 454094 627432
rect 454194 627332 454318 627432
rect 454418 627332 454542 627432
rect 454642 627332 454766 627432
rect 454866 627332 454990 627432
rect 455090 627332 455214 627432
rect 455314 627332 455438 627432
rect 455538 627332 455662 627432
rect 455762 627332 455886 627432
rect 455986 627332 456010 627432
rect 449350 627208 456010 627332
rect 449350 627108 449390 627208
rect 449490 627108 449614 627208
rect 449714 627108 449838 627208
rect 449938 627108 450062 627208
rect 450162 627108 450286 627208
rect 450386 627108 450510 627208
rect 450610 627108 450734 627208
rect 450834 627108 450958 627208
rect 451058 627108 451182 627208
rect 451282 627108 451406 627208
rect 451506 627108 451630 627208
rect 451730 627108 451854 627208
rect 451954 627108 452078 627208
rect 452178 627108 452302 627208
rect 452402 627108 452526 627208
rect 452626 627108 452750 627208
rect 452850 627108 452974 627208
rect 453074 627108 453198 627208
rect 453298 627108 453422 627208
rect 453522 627108 453646 627208
rect 453746 627108 453870 627208
rect 453970 627108 454094 627208
rect 454194 627108 454318 627208
rect 454418 627108 454542 627208
rect 454642 627108 454766 627208
rect 454866 627108 454990 627208
rect 455090 627108 455214 627208
rect 455314 627108 455438 627208
rect 455538 627108 455662 627208
rect 455762 627108 455886 627208
rect 455986 627108 456010 627208
rect 449350 626984 456010 627108
rect 449350 626884 449390 626984
rect 449490 626884 449614 626984
rect 449714 626884 449838 626984
rect 449938 626884 450062 626984
rect 450162 626884 450286 626984
rect 450386 626884 450510 626984
rect 450610 626884 450734 626984
rect 450834 626884 450958 626984
rect 451058 626884 451182 626984
rect 451282 626884 451406 626984
rect 451506 626884 451630 626984
rect 451730 626884 451854 626984
rect 451954 626884 452078 626984
rect 452178 626884 452302 626984
rect 452402 626884 452526 626984
rect 452626 626884 452750 626984
rect 452850 626884 452974 626984
rect 453074 626884 453198 626984
rect 453298 626884 453422 626984
rect 453522 626884 453646 626984
rect 453746 626884 453870 626984
rect 453970 626884 454094 626984
rect 454194 626884 454318 626984
rect 454418 626884 454542 626984
rect 454642 626884 454766 626984
rect 454866 626884 454990 626984
rect 455090 626884 455214 626984
rect 455314 626884 455438 626984
rect 455538 626884 455662 626984
rect 455762 626884 455886 626984
rect 455986 626884 456010 626984
rect 449350 626760 456010 626884
rect 449350 626660 449390 626760
rect 449490 626660 449614 626760
rect 449714 626660 449838 626760
rect 449938 626660 450062 626760
rect 450162 626660 450286 626760
rect 450386 626660 450510 626760
rect 450610 626660 450734 626760
rect 450834 626660 450958 626760
rect 451058 626660 451182 626760
rect 451282 626660 451406 626760
rect 451506 626660 451630 626760
rect 451730 626660 451854 626760
rect 451954 626660 452078 626760
rect 452178 626660 452302 626760
rect 452402 626660 452526 626760
rect 452626 626660 452750 626760
rect 452850 626660 452974 626760
rect 453074 626660 453198 626760
rect 453298 626660 453422 626760
rect 453522 626660 453646 626760
rect 453746 626660 453870 626760
rect 453970 626660 454094 626760
rect 454194 626660 454318 626760
rect 454418 626660 454542 626760
rect 454642 626660 454766 626760
rect 454866 626660 454990 626760
rect 455090 626660 455214 626760
rect 455314 626660 455438 626760
rect 455538 626660 455662 626760
rect 455762 626660 455886 626760
rect 455986 626660 456010 626760
rect 449350 626626 456010 626660
rect 475620 627676 482280 627706
rect 475620 627576 475660 627676
rect 475760 627576 475884 627676
rect 475984 627576 476108 627676
rect 476208 627576 476332 627676
rect 476432 627576 476556 627676
rect 476656 627576 476780 627676
rect 476880 627576 477004 627676
rect 477104 627576 477228 627676
rect 477328 627576 477452 627676
rect 477552 627576 477676 627676
rect 477776 627576 477900 627676
rect 478000 627576 478124 627676
rect 478224 627576 478348 627676
rect 478448 627576 478572 627676
rect 478672 627576 478796 627676
rect 478896 627576 479020 627676
rect 479120 627576 479244 627676
rect 479344 627576 479468 627676
rect 479568 627576 479692 627676
rect 479792 627576 479916 627676
rect 480016 627576 480140 627676
rect 480240 627576 480364 627676
rect 480464 627576 480588 627676
rect 480688 627576 480812 627676
rect 480912 627576 481036 627676
rect 481136 627576 481260 627676
rect 481360 627576 481484 627676
rect 481584 627576 481708 627676
rect 481808 627576 481932 627676
rect 482032 627576 482156 627676
rect 482256 627576 482280 627676
rect 475620 627452 482280 627576
rect 475620 627352 475660 627452
rect 475760 627352 475884 627452
rect 475984 627352 476108 627452
rect 476208 627352 476332 627452
rect 476432 627352 476556 627452
rect 476656 627352 476780 627452
rect 476880 627352 477004 627452
rect 477104 627352 477228 627452
rect 477328 627352 477452 627452
rect 477552 627352 477676 627452
rect 477776 627352 477900 627452
rect 478000 627352 478124 627452
rect 478224 627352 478348 627452
rect 478448 627352 478572 627452
rect 478672 627352 478796 627452
rect 478896 627352 479020 627452
rect 479120 627352 479244 627452
rect 479344 627352 479468 627452
rect 479568 627352 479692 627452
rect 479792 627352 479916 627452
rect 480016 627352 480140 627452
rect 480240 627352 480364 627452
rect 480464 627352 480588 627452
rect 480688 627352 480812 627452
rect 480912 627352 481036 627452
rect 481136 627352 481260 627452
rect 481360 627352 481484 627452
rect 481584 627352 481708 627452
rect 481808 627352 481932 627452
rect 482032 627352 482156 627452
rect 482256 627352 482280 627452
rect 475620 627228 482280 627352
rect 475620 627128 475660 627228
rect 475760 627128 475884 627228
rect 475984 627128 476108 627228
rect 476208 627128 476332 627228
rect 476432 627128 476556 627228
rect 476656 627128 476780 627228
rect 476880 627128 477004 627228
rect 477104 627128 477228 627228
rect 477328 627128 477452 627228
rect 477552 627128 477676 627228
rect 477776 627128 477900 627228
rect 478000 627128 478124 627228
rect 478224 627128 478348 627228
rect 478448 627128 478572 627228
rect 478672 627128 478796 627228
rect 478896 627128 479020 627228
rect 479120 627128 479244 627228
rect 479344 627128 479468 627228
rect 479568 627128 479692 627228
rect 479792 627128 479916 627228
rect 480016 627128 480140 627228
rect 480240 627128 480364 627228
rect 480464 627128 480588 627228
rect 480688 627128 480812 627228
rect 480912 627128 481036 627228
rect 481136 627128 481260 627228
rect 481360 627128 481484 627228
rect 481584 627128 481708 627228
rect 481808 627128 481932 627228
rect 482032 627128 482156 627228
rect 482256 627128 482280 627228
rect 475620 627004 482280 627128
rect 475620 626904 475660 627004
rect 475760 626904 475884 627004
rect 475984 626904 476108 627004
rect 476208 626904 476332 627004
rect 476432 626904 476556 627004
rect 476656 626904 476780 627004
rect 476880 626904 477004 627004
rect 477104 626904 477228 627004
rect 477328 626904 477452 627004
rect 477552 626904 477676 627004
rect 477776 626904 477900 627004
rect 478000 626904 478124 627004
rect 478224 626904 478348 627004
rect 478448 626904 478572 627004
rect 478672 626904 478796 627004
rect 478896 626904 479020 627004
rect 479120 626904 479244 627004
rect 479344 626904 479468 627004
rect 479568 626904 479692 627004
rect 479792 626904 479916 627004
rect 480016 626904 480140 627004
rect 480240 626904 480364 627004
rect 480464 626904 480588 627004
rect 480688 626904 480812 627004
rect 480912 626904 481036 627004
rect 481136 626904 481260 627004
rect 481360 626904 481484 627004
rect 481584 626904 481708 627004
rect 481808 626904 481932 627004
rect 482032 626904 482156 627004
rect 482256 626904 482280 627004
rect 475620 626780 482280 626904
rect 475620 626680 475660 626780
rect 475760 626680 475884 626780
rect 475984 626680 476108 626780
rect 476208 626680 476332 626780
rect 476432 626680 476556 626780
rect 476656 626680 476780 626780
rect 476880 626680 477004 626780
rect 477104 626680 477228 626780
rect 477328 626680 477452 626780
rect 477552 626680 477676 626780
rect 477776 626680 477900 626780
rect 478000 626680 478124 626780
rect 478224 626680 478348 626780
rect 478448 626680 478572 626780
rect 478672 626680 478796 626780
rect 478896 626680 479020 626780
rect 479120 626680 479244 626780
rect 479344 626680 479468 626780
rect 479568 626680 479692 626780
rect 479792 626680 479916 626780
rect 480016 626680 480140 626780
rect 480240 626680 480364 626780
rect 480464 626680 480588 626780
rect 480688 626680 480812 626780
rect 480912 626680 481036 626780
rect 481136 626680 481260 626780
rect 481360 626680 481484 626780
rect 481584 626680 481708 626780
rect 481808 626680 481932 626780
rect 482032 626680 482156 626780
rect 482256 626680 482280 626780
rect 475620 626646 482280 626680
<< via1 >>
rect 438920 654776 439020 654876
rect 439144 654776 439244 654876
rect 439368 654776 439468 654876
rect 439592 654776 439692 654876
rect 439816 654776 439916 654876
rect 440040 654776 440140 654876
rect 440264 654776 440364 654876
rect 440488 654776 440588 654876
rect 440712 654776 440812 654876
rect 440936 654776 441036 654876
rect 441160 654776 441260 654876
rect 441384 654776 441484 654876
rect 441608 654776 441708 654876
rect 441832 654776 441932 654876
rect 442056 654776 442156 654876
rect 442280 654776 442380 654876
rect 442504 654776 442604 654876
rect 442728 654776 442828 654876
rect 442952 654776 443052 654876
rect 443176 654776 443276 654876
rect 443400 654776 443500 654876
rect 443624 654776 443724 654876
rect 443848 654776 443948 654876
rect 444072 654776 444172 654876
rect 444296 654776 444396 654876
rect 444520 654776 444620 654876
rect 444744 654776 444844 654876
rect 444968 654776 445068 654876
rect 445192 654776 445292 654876
rect 445416 654776 445516 654876
rect 438920 654552 439020 654652
rect 439144 654552 439244 654652
rect 439368 654552 439468 654652
rect 439592 654552 439692 654652
rect 439816 654552 439916 654652
rect 440040 654552 440140 654652
rect 440264 654552 440364 654652
rect 440488 654552 440588 654652
rect 440712 654552 440812 654652
rect 440936 654552 441036 654652
rect 441160 654552 441260 654652
rect 441384 654552 441484 654652
rect 441608 654552 441708 654652
rect 441832 654552 441932 654652
rect 442056 654552 442156 654652
rect 442280 654552 442380 654652
rect 442504 654552 442604 654652
rect 442728 654552 442828 654652
rect 442952 654552 443052 654652
rect 443176 654552 443276 654652
rect 443400 654552 443500 654652
rect 443624 654552 443724 654652
rect 443848 654552 443948 654652
rect 444072 654552 444172 654652
rect 444296 654552 444396 654652
rect 444520 654552 444620 654652
rect 444744 654552 444844 654652
rect 444968 654552 445068 654652
rect 445192 654552 445292 654652
rect 445416 654552 445516 654652
rect 438920 654328 439020 654428
rect 439144 654328 439244 654428
rect 439368 654328 439468 654428
rect 439592 654328 439692 654428
rect 439816 654328 439916 654428
rect 440040 654328 440140 654428
rect 440264 654328 440364 654428
rect 440488 654328 440588 654428
rect 440712 654328 440812 654428
rect 440936 654328 441036 654428
rect 441160 654328 441260 654428
rect 441384 654328 441484 654428
rect 441608 654328 441708 654428
rect 441832 654328 441932 654428
rect 442056 654328 442156 654428
rect 442280 654328 442380 654428
rect 442504 654328 442604 654428
rect 442728 654328 442828 654428
rect 442952 654328 443052 654428
rect 443176 654328 443276 654428
rect 443400 654328 443500 654428
rect 443624 654328 443724 654428
rect 443848 654328 443948 654428
rect 444072 654328 444172 654428
rect 444296 654328 444396 654428
rect 444520 654328 444620 654428
rect 444744 654328 444844 654428
rect 444968 654328 445068 654428
rect 445192 654328 445292 654428
rect 445416 654328 445516 654428
rect 438920 654104 439020 654204
rect 439144 654104 439244 654204
rect 439368 654104 439468 654204
rect 439592 654104 439692 654204
rect 439816 654104 439916 654204
rect 440040 654104 440140 654204
rect 440264 654104 440364 654204
rect 440488 654104 440588 654204
rect 440712 654104 440812 654204
rect 440936 654104 441036 654204
rect 441160 654104 441260 654204
rect 441384 654104 441484 654204
rect 441608 654104 441708 654204
rect 441832 654104 441932 654204
rect 442056 654104 442156 654204
rect 442280 654104 442380 654204
rect 442504 654104 442604 654204
rect 442728 654104 442828 654204
rect 442952 654104 443052 654204
rect 443176 654104 443276 654204
rect 443400 654104 443500 654204
rect 443624 654104 443724 654204
rect 443848 654104 443948 654204
rect 444072 654104 444172 654204
rect 444296 654104 444396 654204
rect 444520 654104 444620 654204
rect 444744 654104 444844 654204
rect 444968 654104 445068 654204
rect 445192 654104 445292 654204
rect 445416 654104 445516 654204
rect 438920 653880 439020 653980
rect 439144 653880 439244 653980
rect 439368 653880 439468 653980
rect 439592 653880 439692 653980
rect 439816 653880 439916 653980
rect 440040 653880 440140 653980
rect 440264 653880 440364 653980
rect 440488 653880 440588 653980
rect 440712 653880 440812 653980
rect 440936 653880 441036 653980
rect 441160 653880 441260 653980
rect 441384 653880 441484 653980
rect 441608 653880 441708 653980
rect 441832 653880 441932 653980
rect 442056 653880 442156 653980
rect 442280 653880 442380 653980
rect 442504 653880 442604 653980
rect 442728 653880 442828 653980
rect 442952 653880 443052 653980
rect 443176 653880 443276 653980
rect 443400 653880 443500 653980
rect 443624 653880 443724 653980
rect 443848 653880 443948 653980
rect 444072 653880 444172 653980
rect 444296 653880 444396 653980
rect 444520 653880 444620 653980
rect 444744 653880 444844 653980
rect 444968 653880 445068 653980
rect 445192 653880 445292 653980
rect 445416 653880 445516 653980
rect 449390 654776 449490 654876
rect 449614 654776 449714 654876
rect 449838 654776 449938 654876
rect 450062 654776 450162 654876
rect 450286 654776 450386 654876
rect 450510 654776 450610 654876
rect 450734 654776 450834 654876
rect 450958 654776 451058 654876
rect 451182 654776 451282 654876
rect 451406 654776 451506 654876
rect 451630 654776 451730 654876
rect 451854 654776 451954 654876
rect 452078 654776 452178 654876
rect 452302 654776 452402 654876
rect 452526 654776 452626 654876
rect 452750 654776 452850 654876
rect 452974 654776 453074 654876
rect 453198 654776 453298 654876
rect 453422 654776 453522 654876
rect 453646 654776 453746 654876
rect 453870 654776 453970 654876
rect 454094 654776 454194 654876
rect 454318 654776 454418 654876
rect 454542 654776 454642 654876
rect 454766 654776 454866 654876
rect 454990 654776 455090 654876
rect 455214 654776 455314 654876
rect 455438 654776 455538 654876
rect 455662 654776 455762 654876
rect 455886 654776 455986 654876
rect 449390 654552 449490 654652
rect 449614 654552 449714 654652
rect 449838 654552 449938 654652
rect 450062 654552 450162 654652
rect 450286 654552 450386 654652
rect 450510 654552 450610 654652
rect 450734 654552 450834 654652
rect 450958 654552 451058 654652
rect 451182 654552 451282 654652
rect 451406 654552 451506 654652
rect 451630 654552 451730 654652
rect 451854 654552 451954 654652
rect 452078 654552 452178 654652
rect 452302 654552 452402 654652
rect 452526 654552 452626 654652
rect 452750 654552 452850 654652
rect 452974 654552 453074 654652
rect 453198 654552 453298 654652
rect 453422 654552 453522 654652
rect 453646 654552 453746 654652
rect 453870 654552 453970 654652
rect 454094 654552 454194 654652
rect 454318 654552 454418 654652
rect 454542 654552 454642 654652
rect 454766 654552 454866 654652
rect 454990 654552 455090 654652
rect 455214 654552 455314 654652
rect 455438 654552 455538 654652
rect 455662 654552 455762 654652
rect 455886 654552 455986 654652
rect 449390 654328 449490 654428
rect 449614 654328 449714 654428
rect 449838 654328 449938 654428
rect 450062 654328 450162 654428
rect 450286 654328 450386 654428
rect 450510 654328 450610 654428
rect 450734 654328 450834 654428
rect 450958 654328 451058 654428
rect 451182 654328 451282 654428
rect 451406 654328 451506 654428
rect 451630 654328 451730 654428
rect 451854 654328 451954 654428
rect 452078 654328 452178 654428
rect 452302 654328 452402 654428
rect 452526 654328 452626 654428
rect 452750 654328 452850 654428
rect 452974 654328 453074 654428
rect 453198 654328 453298 654428
rect 453422 654328 453522 654428
rect 453646 654328 453746 654428
rect 453870 654328 453970 654428
rect 454094 654328 454194 654428
rect 454318 654328 454418 654428
rect 454542 654328 454642 654428
rect 454766 654328 454866 654428
rect 454990 654328 455090 654428
rect 455214 654328 455314 654428
rect 455438 654328 455538 654428
rect 455662 654328 455762 654428
rect 455886 654328 455986 654428
rect 449390 654104 449490 654204
rect 449614 654104 449714 654204
rect 449838 654104 449938 654204
rect 450062 654104 450162 654204
rect 450286 654104 450386 654204
rect 450510 654104 450610 654204
rect 450734 654104 450834 654204
rect 450958 654104 451058 654204
rect 451182 654104 451282 654204
rect 451406 654104 451506 654204
rect 451630 654104 451730 654204
rect 451854 654104 451954 654204
rect 452078 654104 452178 654204
rect 452302 654104 452402 654204
rect 452526 654104 452626 654204
rect 452750 654104 452850 654204
rect 452974 654104 453074 654204
rect 453198 654104 453298 654204
rect 453422 654104 453522 654204
rect 453646 654104 453746 654204
rect 453870 654104 453970 654204
rect 454094 654104 454194 654204
rect 454318 654104 454418 654204
rect 454542 654104 454642 654204
rect 454766 654104 454866 654204
rect 454990 654104 455090 654204
rect 455214 654104 455314 654204
rect 455438 654104 455538 654204
rect 455662 654104 455762 654204
rect 455886 654104 455986 654204
rect 449390 653880 449490 653980
rect 449614 653880 449714 653980
rect 449838 653880 449938 653980
rect 450062 653880 450162 653980
rect 450286 653880 450386 653980
rect 450510 653880 450610 653980
rect 450734 653880 450834 653980
rect 450958 653880 451058 653980
rect 451182 653880 451282 653980
rect 451406 653880 451506 653980
rect 451630 653880 451730 653980
rect 451854 653880 451954 653980
rect 452078 653880 452178 653980
rect 452302 653880 452402 653980
rect 452526 653880 452626 653980
rect 452750 653880 452850 653980
rect 452974 653880 453074 653980
rect 453198 653880 453298 653980
rect 453422 653880 453522 653980
rect 453646 653880 453746 653980
rect 453870 653880 453970 653980
rect 454094 653880 454194 653980
rect 454318 653880 454418 653980
rect 454542 653880 454642 653980
rect 454766 653880 454866 653980
rect 454990 653880 455090 653980
rect 455214 653880 455314 653980
rect 455438 653880 455538 653980
rect 455662 653880 455762 653980
rect 455886 653880 455986 653980
rect 475660 654796 475760 654896
rect 475884 654796 475984 654896
rect 476108 654796 476208 654896
rect 476332 654796 476432 654896
rect 476556 654796 476656 654896
rect 476780 654796 476880 654896
rect 477004 654796 477104 654896
rect 477228 654796 477328 654896
rect 477452 654796 477552 654896
rect 477676 654796 477776 654896
rect 477900 654796 478000 654896
rect 478124 654796 478224 654896
rect 478348 654796 478448 654896
rect 478572 654796 478672 654896
rect 478796 654796 478896 654896
rect 479020 654796 479120 654896
rect 479244 654796 479344 654896
rect 479468 654796 479568 654896
rect 479692 654796 479792 654896
rect 479916 654796 480016 654896
rect 480140 654796 480240 654896
rect 480364 654796 480464 654896
rect 480588 654796 480688 654896
rect 480812 654796 480912 654896
rect 481036 654796 481136 654896
rect 481260 654796 481360 654896
rect 481484 654796 481584 654896
rect 481708 654796 481808 654896
rect 481932 654796 482032 654896
rect 482156 654796 482256 654896
rect 475660 654572 475760 654672
rect 475884 654572 475984 654672
rect 476108 654572 476208 654672
rect 476332 654572 476432 654672
rect 476556 654572 476656 654672
rect 476780 654572 476880 654672
rect 477004 654572 477104 654672
rect 477228 654572 477328 654672
rect 477452 654572 477552 654672
rect 477676 654572 477776 654672
rect 477900 654572 478000 654672
rect 478124 654572 478224 654672
rect 478348 654572 478448 654672
rect 478572 654572 478672 654672
rect 478796 654572 478896 654672
rect 479020 654572 479120 654672
rect 479244 654572 479344 654672
rect 479468 654572 479568 654672
rect 479692 654572 479792 654672
rect 479916 654572 480016 654672
rect 480140 654572 480240 654672
rect 480364 654572 480464 654672
rect 480588 654572 480688 654672
rect 480812 654572 480912 654672
rect 481036 654572 481136 654672
rect 481260 654572 481360 654672
rect 481484 654572 481584 654672
rect 481708 654572 481808 654672
rect 481932 654572 482032 654672
rect 482156 654572 482256 654672
rect 475660 654348 475760 654448
rect 475884 654348 475984 654448
rect 476108 654348 476208 654448
rect 476332 654348 476432 654448
rect 476556 654348 476656 654448
rect 476780 654348 476880 654448
rect 477004 654348 477104 654448
rect 477228 654348 477328 654448
rect 477452 654348 477552 654448
rect 477676 654348 477776 654448
rect 477900 654348 478000 654448
rect 478124 654348 478224 654448
rect 478348 654348 478448 654448
rect 478572 654348 478672 654448
rect 478796 654348 478896 654448
rect 479020 654348 479120 654448
rect 479244 654348 479344 654448
rect 479468 654348 479568 654448
rect 479692 654348 479792 654448
rect 479916 654348 480016 654448
rect 480140 654348 480240 654448
rect 480364 654348 480464 654448
rect 480588 654348 480688 654448
rect 480812 654348 480912 654448
rect 481036 654348 481136 654448
rect 481260 654348 481360 654448
rect 481484 654348 481584 654448
rect 481708 654348 481808 654448
rect 481932 654348 482032 654448
rect 482156 654348 482256 654448
rect 475660 654124 475760 654224
rect 475884 654124 475984 654224
rect 476108 654124 476208 654224
rect 476332 654124 476432 654224
rect 476556 654124 476656 654224
rect 476780 654124 476880 654224
rect 477004 654124 477104 654224
rect 477228 654124 477328 654224
rect 477452 654124 477552 654224
rect 477676 654124 477776 654224
rect 477900 654124 478000 654224
rect 478124 654124 478224 654224
rect 478348 654124 478448 654224
rect 478572 654124 478672 654224
rect 478796 654124 478896 654224
rect 479020 654124 479120 654224
rect 479244 654124 479344 654224
rect 479468 654124 479568 654224
rect 479692 654124 479792 654224
rect 479916 654124 480016 654224
rect 480140 654124 480240 654224
rect 480364 654124 480464 654224
rect 480588 654124 480688 654224
rect 480812 654124 480912 654224
rect 481036 654124 481136 654224
rect 481260 654124 481360 654224
rect 481484 654124 481584 654224
rect 481708 654124 481808 654224
rect 481932 654124 482032 654224
rect 482156 654124 482256 654224
rect 475660 653900 475760 654000
rect 475884 653900 475984 654000
rect 476108 653900 476208 654000
rect 476332 653900 476432 654000
rect 476556 653900 476656 654000
rect 476780 653900 476880 654000
rect 477004 653900 477104 654000
rect 477228 653900 477328 654000
rect 477452 653900 477552 654000
rect 477676 653900 477776 654000
rect 477900 653900 478000 654000
rect 478124 653900 478224 654000
rect 478348 653900 478448 654000
rect 478572 653900 478672 654000
rect 478796 653900 478896 654000
rect 479020 653900 479120 654000
rect 479244 653900 479344 654000
rect 479468 653900 479568 654000
rect 479692 653900 479792 654000
rect 479916 653900 480016 654000
rect 480140 653900 480240 654000
rect 480364 653900 480464 654000
rect 480588 653900 480688 654000
rect 480812 653900 480912 654000
rect 481036 653900 481136 654000
rect 481260 653900 481360 654000
rect 481484 653900 481584 654000
rect 481708 653900 481808 654000
rect 481932 653900 482032 654000
rect 482156 653900 482256 654000
rect 440702 652740 451946 652754
rect 440702 651942 440716 652740
rect 440716 651942 451932 652740
rect 451932 651942 451946 652740
rect 440702 651928 451946 651942
rect 463968 650656 464526 651214
rect 465592 650656 466150 651214
rect 469682 650656 470240 651214
rect 472136 650656 472694 651214
rect 437894 650078 437994 650178
rect 438118 650078 438218 650178
rect 438342 650078 438442 650178
rect 438566 650078 438666 650178
rect 438790 650078 438890 650178
rect 437894 649854 437994 649954
rect 438118 649854 438218 649954
rect 438342 649854 438442 649954
rect 438566 649854 438666 649954
rect 438790 649854 438890 649954
rect 457412 649856 457970 650414
rect 463138 649856 463696 650414
rect 466410 649856 466968 650414
rect 468864 649856 469422 650414
rect 471318 649856 471876 650414
rect 473772 649856 474330 650414
rect 482174 650078 482274 650178
rect 482398 650078 482498 650178
rect 482622 650078 482722 650178
rect 482846 650078 482946 650178
rect 483070 650078 483170 650178
rect 482174 649854 482274 649954
rect 482398 649854 482498 649954
rect 482622 649854 482722 649954
rect 482846 649854 482946 649954
rect 483070 649854 483170 649954
rect 437894 649630 437994 649730
rect 438118 649630 438218 649730
rect 438342 649630 438442 649730
rect 438566 649630 438666 649730
rect 438790 649630 438890 649730
rect 437894 649406 437994 649506
rect 438118 649406 438218 649506
rect 438342 649406 438442 649506
rect 438566 649406 438666 649506
rect 438790 649406 438890 649506
rect 437894 649182 437994 649282
rect 438118 649182 438218 649282
rect 438342 649182 438442 649282
rect 438566 649182 438666 649282
rect 438790 649182 438890 649282
rect 457412 649664 457970 649676
rect 457412 649267 457422 649664
rect 457422 649267 457960 649664
rect 457960 649267 457970 649664
rect 457412 649256 457970 649267
rect 458230 649664 458788 649676
rect 458230 649267 458240 649664
rect 458240 649267 458778 649664
rect 458778 649267 458788 649664
rect 458230 649256 458788 649267
rect 482174 649630 482274 649730
rect 482398 649630 482498 649730
rect 482622 649630 482722 649730
rect 482846 649630 482946 649730
rect 483070 649630 483170 649730
rect 462320 649602 462878 649614
rect 462320 649205 462330 649602
rect 462330 649205 462868 649602
rect 462868 649205 462878 649602
rect 462320 649194 462878 649205
rect 463138 649602 463696 649614
rect 463138 649205 463148 649602
rect 463148 649205 463686 649602
rect 463686 649205 463696 649602
rect 463138 649194 463696 649205
rect 463956 649602 464514 649614
rect 463956 649205 463966 649602
rect 463966 649205 464504 649602
rect 464504 649205 464514 649602
rect 463956 649194 464514 649205
rect 464774 649602 465332 649614
rect 464774 649205 464784 649602
rect 464784 649205 465322 649602
rect 465322 649205 465332 649602
rect 464774 649194 465332 649205
rect 465592 649602 466150 649614
rect 465592 649205 465602 649602
rect 465602 649205 466140 649602
rect 466140 649205 466150 649602
rect 465592 649194 466150 649205
rect 466410 649602 466968 649614
rect 466410 649205 466420 649602
rect 466420 649205 466958 649602
rect 466958 649205 466968 649602
rect 466410 649194 466968 649205
rect 467228 649602 467786 649614
rect 467228 649205 467238 649602
rect 467238 649205 467776 649602
rect 467776 649205 467786 649602
rect 467228 649194 467786 649205
rect 468046 649602 468604 649614
rect 468046 649205 468056 649602
rect 468056 649205 468594 649602
rect 468594 649205 468604 649602
rect 468046 649194 468604 649205
rect 468864 649602 469422 649614
rect 468864 649205 468874 649602
rect 468874 649205 469412 649602
rect 469412 649205 469422 649602
rect 468864 649194 469422 649205
rect 469682 649602 470240 649614
rect 469682 649205 469692 649602
rect 469692 649205 470230 649602
rect 470230 649205 470240 649602
rect 469682 649194 470240 649205
rect 470500 649602 471058 649614
rect 470500 649205 470510 649602
rect 470510 649205 471048 649602
rect 471048 649205 471058 649602
rect 470500 649194 471058 649205
rect 471318 649602 471876 649614
rect 471318 649205 471328 649602
rect 471328 649205 471866 649602
rect 471866 649205 471876 649602
rect 471318 649194 471876 649205
rect 472136 649602 472694 649614
rect 472136 649205 472146 649602
rect 472146 649205 472684 649602
rect 472684 649205 472694 649602
rect 472136 649194 472694 649205
rect 472954 649602 473512 649614
rect 472954 649205 472964 649602
rect 472964 649205 473502 649602
rect 473502 649205 473512 649602
rect 472954 649194 473512 649205
rect 473772 649602 474330 649614
rect 473772 649205 473782 649602
rect 473782 649205 474320 649602
rect 474320 649205 474330 649602
rect 473772 649194 474330 649205
rect 482174 649406 482274 649506
rect 482398 649406 482498 649506
rect 482622 649406 482722 649506
rect 482846 649406 482946 649506
rect 483070 649406 483170 649506
rect 437894 648958 437994 649058
rect 438118 648958 438218 649058
rect 438342 648958 438442 649058
rect 438566 648958 438666 649058
rect 438790 648958 438890 649058
rect 482174 649182 482274 649282
rect 482398 649182 482498 649282
rect 482622 649182 482722 649282
rect 482846 649182 482946 649282
rect 483070 649182 483170 649282
rect 482174 648958 482274 649058
rect 482398 648958 482498 649058
rect 482622 648958 482722 649058
rect 482846 648958 482946 649058
rect 483070 648958 483170 649058
rect 437894 648734 437994 648834
rect 438118 648734 438218 648834
rect 438342 648734 438442 648834
rect 438566 648734 438666 648834
rect 438790 648734 438890 648834
rect 437894 648510 437994 648610
rect 438118 648510 438218 648610
rect 438342 648510 438442 648610
rect 438566 648510 438666 648610
rect 438790 648510 438890 648610
rect 458230 648460 458788 648952
rect 462320 648394 462878 648952
rect 464774 648394 465332 648952
rect 467228 648394 467786 648952
rect 470500 648394 471058 648952
rect 472954 648394 473512 648952
rect 482174 648734 482274 648834
rect 482398 648734 482498 648834
rect 482622 648734 482722 648834
rect 482846 648734 482946 648834
rect 483070 648734 483170 648834
rect 482174 648510 482274 648610
rect 482398 648510 482498 648610
rect 482622 648510 482722 648610
rect 482846 648510 482946 648610
rect 483070 648510 483170 648610
rect 437894 648286 437994 648386
rect 438118 648286 438218 648386
rect 438342 648286 438442 648386
rect 438566 648286 438666 648386
rect 438790 648286 438890 648386
rect 482174 648286 482274 648386
rect 482398 648286 482498 648386
rect 482622 648286 482722 648386
rect 482846 648286 482946 648386
rect 483070 648286 483170 648386
rect 437894 648062 437994 648162
rect 438118 648062 438218 648162
rect 438342 648062 438442 648162
rect 438566 648062 438666 648162
rect 438790 648062 438890 648162
rect 437894 647838 437994 647938
rect 438118 647838 438218 647938
rect 438342 647838 438442 647938
rect 438566 647838 438666 647938
rect 438790 647838 438890 647938
rect 482174 648062 482274 648162
rect 482398 648062 482498 648162
rect 482622 648062 482722 648162
rect 482846 648062 482946 648162
rect 483070 648062 483170 648162
rect 437894 647614 437994 647714
rect 438118 647614 438218 647714
rect 438342 647614 438442 647714
rect 438566 647614 438666 647714
rect 438790 647614 438890 647714
rect 437894 647390 437994 647490
rect 438118 647390 438218 647490
rect 438342 647390 438442 647490
rect 438566 647390 438666 647490
rect 438790 647390 438890 647490
rect 437894 647166 437994 647266
rect 438118 647166 438218 647266
rect 438342 647166 438442 647266
rect 438566 647166 438666 647266
rect 438790 647166 438890 647266
rect 437894 646942 437994 647042
rect 438118 646942 438218 647042
rect 438342 646942 438442 647042
rect 438566 646942 438666 647042
rect 438790 646942 438890 647042
rect 437894 646718 437994 646818
rect 438118 646718 438218 646818
rect 438342 646718 438442 646818
rect 438566 646718 438666 646818
rect 438790 646718 438890 646818
rect 437894 646494 437994 646594
rect 438118 646494 438218 646594
rect 438342 646494 438442 646594
rect 438566 646494 438666 646594
rect 438790 646494 438890 646594
rect 437894 646270 437994 646370
rect 438118 646270 438218 646370
rect 438342 646270 438442 646370
rect 438566 646270 438666 646370
rect 438790 646270 438890 646370
rect 437894 646046 437994 646146
rect 438118 646046 438218 646146
rect 438342 646046 438442 646146
rect 438566 646046 438666 646146
rect 438790 646046 438890 646146
rect 437894 645822 437994 645922
rect 438118 645822 438218 645922
rect 438342 645822 438442 645922
rect 438566 645822 438666 645922
rect 438790 645822 438890 645922
rect 437894 645598 437994 645698
rect 438118 645598 438218 645698
rect 438342 645598 438442 645698
rect 438566 645598 438666 645698
rect 438790 645598 438890 645698
rect 437894 645374 437994 645474
rect 438118 645374 438218 645474
rect 438342 645374 438442 645474
rect 438566 645374 438666 645474
rect 438790 645374 438890 645474
rect 437894 645150 437994 645250
rect 438118 645150 438218 645250
rect 438342 645150 438442 645250
rect 438566 645150 438666 645250
rect 438790 645150 438890 645250
rect 437894 644926 437994 645026
rect 438118 644926 438218 645026
rect 438342 644926 438442 645026
rect 438566 644926 438666 645026
rect 438790 644926 438890 645026
rect 482174 647838 482274 647938
rect 482398 647838 482498 647938
rect 482622 647838 482722 647938
rect 482846 647838 482946 647938
rect 483070 647838 483170 647938
rect 482174 647614 482274 647714
rect 482398 647614 482498 647714
rect 482622 647614 482722 647714
rect 482846 647614 482946 647714
rect 483070 647614 483170 647714
rect 482174 647390 482274 647490
rect 482398 647390 482498 647490
rect 482622 647390 482722 647490
rect 482846 647390 482946 647490
rect 483070 647390 483170 647490
rect 482174 647166 482274 647266
rect 482398 647166 482498 647266
rect 482622 647166 482722 647266
rect 482846 647166 482946 647266
rect 483070 647166 483170 647266
rect 482174 646942 482274 647042
rect 482398 646942 482498 647042
rect 482622 646942 482722 647042
rect 482846 646942 482946 647042
rect 483070 646942 483170 647042
rect 482174 646718 482274 646818
rect 482398 646718 482498 646818
rect 482622 646718 482722 646818
rect 482846 646718 482946 646818
rect 483070 646718 483170 646818
rect 482174 646494 482274 646594
rect 482398 646494 482498 646594
rect 482622 646494 482722 646594
rect 482846 646494 482946 646594
rect 483070 646494 483170 646594
rect 482174 646270 482274 646370
rect 482398 646270 482498 646370
rect 482622 646270 482722 646370
rect 482846 646270 482946 646370
rect 483070 646270 483170 646370
rect 482174 646046 482274 646146
rect 482398 646046 482498 646146
rect 482622 646046 482722 646146
rect 482846 646046 482946 646146
rect 483070 646046 483170 646146
rect 482174 645822 482274 645922
rect 482398 645822 482498 645922
rect 482622 645822 482722 645922
rect 482846 645822 482946 645922
rect 483070 645822 483170 645922
rect 482174 645598 482274 645698
rect 482398 645598 482498 645698
rect 482622 645598 482722 645698
rect 482846 645598 482946 645698
rect 483070 645598 483170 645698
rect 482174 645374 482274 645474
rect 482398 645374 482498 645474
rect 482622 645374 482722 645474
rect 482846 645374 482946 645474
rect 483070 645374 483170 645474
rect 482174 645150 482274 645250
rect 482398 645150 482498 645250
rect 482622 645150 482722 645250
rect 482846 645150 482946 645250
rect 483070 645150 483170 645250
rect 437894 644702 437994 644802
rect 438118 644702 438218 644802
rect 438342 644702 438442 644802
rect 438566 644702 438666 644802
rect 438790 644702 438890 644802
rect 437894 644478 437994 644578
rect 438118 644478 438218 644578
rect 438342 644478 438442 644578
rect 438566 644478 438666 644578
rect 438790 644478 438890 644578
rect 437894 644254 437994 644354
rect 438118 644254 438218 644354
rect 438342 644254 438442 644354
rect 438566 644254 438666 644354
rect 438790 644254 438890 644354
rect 437894 644030 437994 644130
rect 438118 644030 438218 644130
rect 438342 644030 438442 644130
rect 438566 644030 438666 644130
rect 438790 644030 438890 644130
rect 437894 643806 437994 643906
rect 438118 643806 438218 643906
rect 438342 643806 438442 643906
rect 438566 643806 438666 643906
rect 438790 643806 438890 643906
rect 437894 643582 437994 643682
rect 438118 643582 438218 643682
rect 438342 643582 438442 643682
rect 438566 643582 438666 643682
rect 438790 643582 438890 643682
rect 482174 644926 482274 645026
rect 482398 644926 482498 645026
rect 482622 644926 482722 645026
rect 482846 644926 482946 645026
rect 483070 644926 483170 645026
rect 482174 644702 482274 644802
rect 482398 644702 482498 644802
rect 482622 644702 482722 644802
rect 482846 644702 482946 644802
rect 483070 644702 483170 644802
rect 463138 643920 463696 644478
rect 466410 643920 466968 644478
rect 468864 643920 469422 644478
rect 471318 643920 471876 644478
rect 482174 644478 482274 644578
rect 482398 644478 482498 644578
rect 482622 644478 482722 644578
rect 482846 644478 482946 644578
rect 483070 644478 483170 644578
rect 482174 644254 482274 644354
rect 482398 644254 482498 644354
rect 482622 644254 482722 644354
rect 482846 644254 482946 644354
rect 483070 644254 483170 644354
rect 482174 644030 482274 644130
rect 482398 644030 482498 644130
rect 482622 644030 482722 644130
rect 482846 644030 482946 644130
rect 483070 644030 483170 644130
rect 482174 643806 482274 643906
rect 482398 643806 482498 643906
rect 482622 643806 482722 643906
rect 482846 643806 482946 643906
rect 483070 643806 483170 643906
rect 463956 643120 464514 643678
rect 465592 643120 466150 643678
rect 469682 643120 470240 643678
rect 482174 643582 482274 643682
rect 482398 643582 482498 643682
rect 482622 643582 482722 643682
rect 482846 643582 482946 643682
rect 483070 643582 483170 643682
rect 462320 642867 462878 642878
rect 462320 642469 462330 642867
rect 462330 642469 462868 642867
rect 462868 642469 462878 642867
rect 462320 642458 462878 642469
rect 463138 642867 463696 642878
rect 463138 642470 463148 642867
rect 463148 642470 463686 642867
rect 463686 642470 463696 642867
rect 463138 642458 463696 642470
rect 463956 642867 464514 642878
rect 463956 642470 463966 642867
rect 463966 642470 464504 642867
rect 464504 642470 464514 642867
rect 463956 642458 464514 642470
rect 464774 642867 465332 642878
rect 464774 642469 464784 642867
rect 464784 642469 465322 642867
rect 465322 642469 465332 642867
rect 464774 642458 465332 642469
rect 465592 642867 466150 642878
rect 465592 642470 465602 642867
rect 465602 642470 466140 642867
rect 466140 642470 466150 642867
rect 465592 642458 466150 642470
rect 466410 642867 466968 642878
rect 466410 642470 466420 642867
rect 466420 642470 466958 642867
rect 466958 642470 466968 642867
rect 466410 642458 466968 642470
rect 467228 642867 467786 642878
rect 467228 642469 467238 642867
rect 467238 642469 467776 642867
rect 467776 642469 467786 642867
rect 467228 642458 467786 642469
rect 468046 642867 468604 642878
rect 468046 642846 468056 642867
rect 467968 642470 468056 642846
rect 468056 642470 468594 642867
rect 468594 642846 468604 642867
rect 468594 642470 468660 642846
rect 467968 642328 468660 642470
rect 468864 642867 469422 642878
rect 468864 642470 468874 642867
rect 468874 642470 469412 642867
rect 469412 642470 469422 642867
rect 468864 642458 469422 642470
rect 469682 642867 470240 642878
rect 469682 642470 469692 642867
rect 469692 642470 470230 642867
rect 470230 642470 470240 642867
rect 469682 642458 470240 642470
rect 470500 642867 471058 642878
rect 470500 642469 470510 642867
rect 470510 642469 471048 642867
rect 471048 642469 471058 642867
rect 470500 642458 471058 642469
rect 471318 642867 471876 642878
rect 471318 642470 471328 642867
rect 471328 642470 471866 642867
rect 471866 642470 471876 642867
rect 471318 642458 471876 642470
rect 462320 641658 462878 642216
rect 464774 641658 465332 642216
rect 467228 641658 467786 642216
rect 470500 641658 471058 642216
rect 472058 642867 472750 642878
rect 472058 642470 472146 642867
rect 472146 642470 472684 642867
rect 472684 642470 472750 642867
rect 472058 642186 472750 642470
rect 459444 640850 459644 641050
rect 459878 640850 460078 641050
rect 460312 640850 460512 641050
rect 460746 640850 460946 641050
rect 461180 640850 461380 641050
rect 461614 640850 461814 641050
rect 462048 640850 462248 641050
rect 462482 640850 462682 641050
rect 462916 640850 463116 641050
rect 463350 640850 463550 641050
rect 463784 640850 463984 641050
rect 464184 640850 464384 641050
rect 464584 640850 464784 641050
rect 464984 640850 465184 641050
rect 465384 640850 465584 641050
rect 465784 640850 465984 641050
rect 466184 640850 466384 641050
rect 466584 640850 466784 641050
rect 466984 640850 467184 641050
rect 467384 640850 467584 641050
rect 468984 640850 469184 641050
rect 469384 640850 469584 641050
rect 469784 640850 469984 641050
rect 470184 640850 470384 641050
rect 470584 640850 470784 641050
rect 470984 640850 471184 641050
rect 471384 640850 471584 641050
rect 471784 640850 471984 641050
rect 472184 640850 472384 641050
rect 459444 640416 459644 640616
rect 459878 640416 460078 640616
rect 460312 640416 460512 640616
rect 460746 640416 460946 640616
rect 461180 640416 461380 640616
rect 461614 640416 461814 640616
rect 462048 640416 462248 640616
rect 462482 640416 462682 640616
rect 462916 640416 463116 640616
rect 463350 640416 463550 640616
rect 463784 640416 463984 640616
rect 472876 642867 473568 642878
rect 472876 642470 472964 642867
rect 472964 642470 473502 642867
rect 473502 642470 473568 642867
rect 472876 642186 473568 642470
rect 459444 639982 459644 640182
rect 459878 639982 460078 640182
rect 460312 639982 460512 640182
rect 460746 639982 460946 640182
rect 461180 639982 461380 640182
rect 461614 639982 461814 640182
rect 462048 639982 462248 640182
rect 462482 639982 462682 640182
rect 462916 639982 463116 640182
rect 463350 639982 463550 640182
rect 463784 639982 463984 640182
rect 453864 639098 455852 639548
rect 452346 638378 452466 638792
rect 451890 637794 452010 638086
rect 437894 636678 437994 636778
rect 438118 636678 438218 636778
rect 438342 636678 438442 636778
rect 438566 636678 438666 636778
rect 438790 636678 438890 636778
rect 437894 636454 437994 636554
rect 438118 636454 438218 636554
rect 438342 636454 438442 636554
rect 438566 636454 438666 636554
rect 438790 636454 438890 636554
rect 437894 636230 437994 636330
rect 438118 636230 438218 636330
rect 438342 636230 438442 636330
rect 438566 636230 438666 636330
rect 438790 636230 438890 636330
rect 443016 636296 443076 636366
rect 443088 636296 443148 636366
rect 443160 636296 443220 636366
rect 443232 636296 443292 636366
rect 443304 636296 443364 636366
rect 443376 636296 443436 636366
rect 443448 636296 443508 636366
rect 443520 636296 443580 636366
rect 443016 636202 443076 636272
rect 443088 636202 443148 636272
rect 443160 636202 443220 636272
rect 443232 636202 443292 636272
rect 443304 636202 443364 636272
rect 443376 636202 443436 636272
rect 443448 636202 443508 636272
rect 443520 636202 443580 636272
rect 437894 636006 437994 636106
rect 438118 636006 438218 636106
rect 438342 636006 438442 636106
rect 438566 636006 438666 636106
rect 438790 636006 438890 636106
rect 437894 635782 437994 635882
rect 438118 635782 438218 635882
rect 438342 635782 438442 635882
rect 438566 635782 438666 635882
rect 438790 635782 438890 635882
rect 437894 635558 437994 635658
rect 438118 635558 438218 635658
rect 438342 635558 438442 635658
rect 438566 635558 438666 635658
rect 438790 635558 438890 635658
rect 437894 635334 437994 635434
rect 438118 635334 438218 635434
rect 438342 635334 438442 635434
rect 438566 635334 438666 635434
rect 438790 635334 438890 635434
rect 437894 635110 437994 635210
rect 438118 635110 438218 635210
rect 438342 635110 438442 635210
rect 438566 635110 438666 635210
rect 438790 635110 438890 635210
rect 437894 634886 437994 634986
rect 438118 634886 438218 634986
rect 438342 634886 438442 634986
rect 438566 634886 438666 634986
rect 438790 634886 438890 634986
rect 437894 634662 437994 634762
rect 438118 634662 438218 634762
rect 438342 634662 438442 634762
rect 438566 634662 438666 634762
rect 438790 634662 438890 634762
rect 437894 634438 437994 634538
rect 438118 634438 438218 634538
rect 438342 634438 438442 634538
rect 438566 634438 438666 634538
rect 438790 634438 438890 634538
rect 437894 634214 437994 634314
rect 438118 634214 438218 634314
rect 438342 634214 438442 634314
rect 438566 634214 438666 634314
rect 438790 634214 438890 634314
rect 437894 633990 437994 634090
rect 438118 633990 438218 634090
rect 438342 633990 438442 634090
rect 438566 633990 438666 634090
rect 438790 633990 438890 634090
rect 437894 633766 437994 633866
rect 438118 633766 438218 633866
rect 438342 633766 438442 633866
rect 438566 633766 438666 633866
rect 438790 633766 438890 633866
rect 437894 633542 437994 633642
rect 438118 633542 438218 633642
rect 438342 633542 438442 633642
rect 438566 633542 438666 633642
rect 438790 633542 438890 633642
rect 437894 633318 437994 633418
rect 438118 633318 438218 633418
rect 438342 633318 438442 633418
rect 438566 633318 438666 633418
rect 438790 633318 438890 633418
rect 437894 633094 437994 633194
rect 438118 633094 438218 633194
rect 438342 633094 438442 633194
rect 438566 633094 438666 633194
rect 438790 633094 438890 633194
rect 437894 632870 437994 632970
rect 438118 632870 438218 632970
rect 438342 632870 438442 632970
rect 438566 632870 438666 632970
rect 438790 632870 438890 632970
rect 437894 632646 437994 632746
rect 438118 632646 438218 632746
rect 438342 632646 438442 632746
rect 438566 632646 438666 632746
rect 438790 632646 438890 632746
rect 440884 632632 440936 632684
rect 437894 632422 437994 632522
rect 438118 632422 438218 632522
rect 438342 632422 438442 632522
rect 438566 632422 438666 632522
rect 438790 632422 438890 632522
rect 442718 632638 442770 632690
rect 443324 632632 443518 632690
rect 441802 632426 441854 632478
rect 437894 632198 437994 632298
rect 438118 632198 438218 632298
rect 438342 632198 438442 632298
rect 438566 632198 438666 632298
rect 438790 632198 438890 632298
rect 437894 631974 437994 632074
rect 438118 631974 438218 632074
rect 438342 631974 438442 632074
rect 438566 631974 438666 632074
rect 438790 631974 438890 632074
rect 437894 631750 437994 631850
rect 438118 631750 438218 631850
rect 438342 631750 438442 631850
rect 438566 631750 438666 631850
rect 438790 631750 438890 631850
rect 437894 631526 437994 631626
rect 438118 631526 438218 631626
rect 438342 631526 438442 631626
rect 438566 631526 438666 631626
rect 438790 631526 438890 631626
rect 437894 631302 437994 631402
rect 438118 631302 438218 631402
rect 438342 631302 438442 631402
rect 438566 631302 438666 631402
rect 438790 631302 438890 631402
rect 437894 631078 437994 631178
rect 438118 631078 438218 631178
rect 438342 631078 438442 631178
rect 438566 631078 438666 631178
rect 438790 631078 438890 631178
rect 437894 630854 437994 630954
rect 438118 630854 438218 630954
rect 438342 630854 438442 630954
rect 438566 630854 438666 630954
rect 438790 630854 438890 630954
rect 437894 630630 437994 630730
rect 438118 630630 438218 630730
rect 438342 630630 438442 630730
rect 438566 630630 438666 630730
rect 438790 630630 438890 630730
rect 437894 630406 437994 630506
rect 438118 630406 438218 630506
rect 438342 630406 438442 630506
rect 438566 630406 438666 630506
rect 438790 630406 438890 630506
rect 437894 630182 437994 630282
rect 438118 630182 438218 630282
rect 438342 630182 438442 630282
rect 438566 630182 438666 630282
rect 438790 630182 438890 630282
rect 443008 629136 443060 629240
rect 446684 634620 446828 634674
rect 446112 634480 446256 634534
rect 447828 634620 447972 634674
rect 447256 634480 447400 634534
rect 448972 634620 449116 634674
rect 448400 634480 448544 634534
rect 444480 632064 444532 632318
rect 445040 632064 445092 632318
rect 445600 632064 445652 632318
rect 446380 632364 446432 632468
rect 446952 632364 447004 632468
rect 446500 632064 446552 632318
rect 446078 632011 446286 632028
rect 446078 631977 446082 632011
rect 446082 631977 446266 632011
rect 446266 631977 446286 632011
rect 446078 631970 446286 631977
rect 446650 632011 446858 632024
rect 446650 631977 446654 632011
rect 446654 631977 446838 632011
rect 446838 631977 446858 632011
rect 446650 631966 446858 631977
rect 447524 632364 447576 632468
rect 448096 632364 448148 632468
rect 447644 632064 447696 632318
rect 447222 632011 447430 632028
rect 447222 631977 447226 632011
rect 447226 631977 447410 632011
rect 447410 631977 447430 632011
rect 447222 631970 447430 631977
rect 447794 632011 448002 632028
rect 447794 631977 447798 632011
rect 447798 631977 447982 632011
rect 447982 631977 448002 632011
rect 447794 631970 448002 631977
rect 448668 632364 448720 632468
rect 449240 632364 449292 632468
rect 448788 632064 448840 632318
rect 449588 632064 449640 632318
rect 448366 632011 448574 632028
rect 448366 631977 448370 632011
rect 448370 631977 448554 632011
rect 448554 631977 448574 632011
rect 448366 631970 448574 631977
rect 448938 632011 449146 632028
rect 448938 631977 448942 632011
rect 448942 631977 449126 632011
rect 449126 631977 449146 632011
rect 448938 631970 449146 631977
rect 450148 632064 450200 632318
rect 453864 638396 455852 638684
rect 456564 637796 458552 638084
rect 452346 634614 452466 634694
rect 451890 634474 452000 634554
rect 450708 632064 450760 632318
rect 452758 632064 453226 632318
rect 443630 629136 443682 629240
rect 444088 629136 444140 629240
rect 444664 629136 444716 629240
rect 445236 629136 445288 629240
rect 445808 629136 445860 629240
rect 446380 629136 446432 629240
rect 446952 629136 447004 629240
rect 447524 629136 447576 629240
rect 448096 629136 448148 629240
rect 448668 629136 448720 629240
rect 449240 629136 449292 629240
rect 449812 629136 449864 629240
rect 450384 629136 450436 629240
rect 450956 629136 451008 629240
rect 451066 629136 451118 629240
rect 451524 629136 451576 629240
rect 452136 629136 452188 629240
rect 452758 629076 453226 629224
rect 471534 639810 472468 640328
rect 467564 639098 469552 639548
rect 467564 638396 469552 638684
rect 464864 637796 466852 638084
rect 443324 628932 443518 629046
rect 444204 628936 444256 629040
rect 444776 628936 444828 629040
rect 445348 628936 445400 629040
rect 449352 628936 449404 629040
rect 449924 628936 449976 629040
rect 450496 628936 450548 629040
rect 454078 629090 454218 629210
rect 454538 629090 454678 629210
rect 454998 629090 455138 629210
rect 455458 629090 455598 629210
rect 455918 629090 456058 629210
rect 456378 629090 456518 629210
rect 456838 629090 456978 629210
rect 457298 629090 457438 629210
rect 457758 629090 457898 629210
rect 458218 629090 458358 629210
rect 459578 629090 459718 629210
rect 460038 629090 460178 629210
rect 460498 629090 460638 629210
rect 460958 629090 461098 629210
rect 461418 629090 461558 629210
rect 461878 629090 462018 629210
rect 462338 629090 462478 629210
rect 462798 629090 462938 629210
rect 463258 629090 463398 629210
rect 463718 629090 463858 629210
rect 465078 629090 465218 629210
rect 465538 629090 465678 629210
rect 465998 629090 466138 629210
rect 466458 629090 466598 629210
rect 466918 629090 467058 629210
rect 467378 629090 467518 629210
rect 467838 629090 467978 629210
rect 468298 629090 468438 629210
rect 468758 629090 468898 629210
rect 472876 639098 473568 639548
rect 473694 642867 474386 642878
rect 473694 642470 473782 642867
rect 473782 642470 474320 642867
rect 474320 642470 474386 642867
rect 473694 642186 474386 642470
rect 473696 637796 474386 638084
rect 472876 635068 473568 635760
rect 471532 629914 472468 630850
rect 477640 635650 477692 635702
rect 477744 635650 477796 635702
rect 477848 635650 477900 635702
rect 477952 635650 478004 635702
rect 478056 635650 478108 635702
rect 478160 635650 478212 635702
rect 477640 635546 477692 635598
rect 477744 635546 477796 635598
rect 477848 635546 477900 635598
rect 477952 635546 478004 635598
rect 478056 635546 478108 635598
rect 478160 635546 478212 635598
rect 477640 635442 477692 635494
rect 477744 635442 477796 635494
rect 477848 635442 477900 635494
rect 477952 635442 478004 635494
rect 478056 635442 478108 635494
rect 478160 635442 478212 635494
rect 477640 635338 477692 635390
rect 477744 635338 477796 635390
rect 477848 635338 477900 635390
rect 477952 635338 478004 635390
rect 478056 635338 478108 635390
rect 478160 635338 478212 635390
rect 477640 635234 477692 635286
rect 477744 635234 477796 635286
rect 477848 635234 477900 635286
rect 477952 635234 478004 635286
rect 478056 635234 478108 635286
rect 478160 635234 478212 635286
rect 477640 635130 477692 635182
rect 477744 635130 477796 635182
rect 477848 635130 477900 635182
rect 477952 635130 478004 635182
rect 478056 635130 478108 635182
rect 478160 635130 478212 635182
rect 476352 630498 476404 630550
rect 476456 630498 476508 630550
rect 476560 630498 476612 630550
rect 476664 630498 476716 630550
rect 476768 630498 476820 630550
rect 476872 630498 476924 630550
rect 476352 630394 476404 630446
rect 476456 630394 476508 630446
rect 476560 630394 476612 630446
rect 476664 630394 476716 630446
rect 476768 630394 476820 630446
rect 476872 630394 476924 630446
rect 476352 630290 476404 630342
rect 476456 630290 476508 630342
rect 476560 630290 476612 630342
rect 476664 630290 476716 630342
rect 476768 630290 476820 630342
rect 476872 630290 476924 630342
rect 476352 630186 476404 630238
rect 476456 630186 476508 630238
rect 476560 630186 476612 630238
rect 476664 630186 476716 630238
rect 476768 630186 476820 630238
rect 476872 630186 476924 630238
rect 482174 636678 482274 636778
rect 482398 636678 482498 636778
rect 482622 636678 482722 636778
rect 482846 636678 482946 636778
rect 483070 636678 483170 636778
rect 482174 636454 482274 636554
rect 482398 636454 482498 636554
rect 482622 636454 482722 636554
rect 482846 636454 482946 636554
rect 483070 636454 483170 636554
rect 482174 636230 482274 636330
rect 482398 636230 482498 636330
rect 482622 636230 482722 636330
rect 482846 636230 482946 636330
rect 483070 636230 483170 636330
rect 482174 636006 482274 636106
rect 482398 636006 482498 636106
rect 482622 636006 482722 636106
rect 482846 636006 482946 636106
rect 483070 636006 483170 636106
rect 482174 635782 482274 635882
rect 482398 635782 482498 635882
rect 482622 635782 482722 635882
rect 482846 635782 482946 635882
rect 483070 635782 483170 635882
rect 482174 635558 482274 635658
rect 482398 635558 482498 635658
rect 482622 635558 482722 635658
rect 482846 635558 482946 635658
rect 483070 635558 483170 635658
rect 482174 635334 482274 635434
rect 482398 635334 482498 635434
rect 482622 635334 482722 635434
rect 482846 635334 482946 635434
rect 483070 635334 483170 635434
rect 482174 635110 482274 635210
rect 482398 635110 482498 635210
rect 482622 635110 482722 635210
rect 482846 635110 482946 635210
rect 483070 635110 483170 635210
rect 482174 634886 482274 634986
rect 482398 634886 482498 634986
rect 482622 634886 482722 634986
rect 482846 634886 482946 634986
rect 483070 634886 483170 634986
rect 482174 634662 482274 634762
rect 482398 634662 482498 634762
rect 482622 634662 482722 634762
rect 482846 634662 482946 634762
rect 483070 634662 483170 634762
rect 482174 634438 482274 634538
rect 482398 634438 482498 634538
rect 482622 634438 482722 634538
rect 482846 634438 482946 634538
rect 483070 634438 483170 634538
rect 482174 634214 482274 634314
rect 482398 634214 482498 634314
rect 482622 634214 482722 634314
rect 482846 634214 482946 634314
rect 483070 634214 483170 634314
rect 482174 633990 482274 634090
rect 482398 633990 482498 634090
rect 482622 633990 482722 634090
rect 482846 633990 482946 634090
rect 483070 633990 483170 634090
rect 482174 633766 482274 633866
rect 482398 633766 482498 633866
rect 482622 633766 482722 633866
rect 482846 633766 482946 633866
rect 483070 633766 483170 633866
rect 482174 633542 482274 633642
rect 482398 633542 482498 633642
rect 482622 633542 482722 633642
rect 482846 633542 482946 633642
rect 483070 633542 483170 633642
rect 482174 633318 482274 633418
rect 482398 633318 482498 633418
rect 482622 633318 482722 633418
rect 482846 633318 482946 633418
rect 483070 633318 483170 633418
rect 482174 633094 482274 633194
rect 482398 633094 482498 633194
rect 482622 633094 482722 633194
rect 482846 633094 482946 633194
rect 483070 633094 483170 633194
rect 482174 632870 482274 632970
rect 482398 632870 482498 632970
rect 482622 632870 482722 632970
rect 482846 632870 482946 632970
rect 483070 632870 483170 632970
rect 482174 632646 482274 632746
rect 482398 632646 482498 632746
rect 482622 632646 482722 632746
rect 482846 632646 482946 632746
rect 483070 632646 483170 632746
rect 482174 632422 482274 632522
rect 482398 632422 482498 632522
rect 482622 632422 482722 632522
rect 482846 632422 482946 632522
rect 483070 632422 483170 632522
rect 482174 632198 482274 632298
rect 482398 632198 482498 632298
rect 482622 632198 482722 632298
rect 482846 632198 482946 632298
rect 483070 632198 483170 632298
rect 482174 631974 482274 632074
rect 482398 631974 482498 632074
rect 482622 631974 482722 632074
rect 482846 631974 482946 632074
rect 483070 631974 483170 632074
rect 482174 631750 482274 631850
rect 482398 631750 482498 631850
rect 482622 631750 482722 631850
rect 482846 631750 482946 631850
rect 483070 631750 483170 631850
rect 482174 631526 482274 631626
rect 482398 631526 482498 631626
rect 482622 631526 482722 631626
rect 482846 631526 482946 631626
rect 483070 631526 483170 631626
rect 482174 631302 482274 631402
rect 482398 631302 482498 631402
rect 482622 631302 482722 631402
rect 482846 631302 482946 631402
rect 483070 631302 483170 631402
rect 482174 631078 482274 631178
rect 482398 631078 482498 631178
rect 482622 631078 482722 631178
rect 482846 631078 482946 631178
rect 483070 631078 483170 631178
rect 482174 630854 482274 630954
rect 482398 630854 482498 630954
rect 482622 630854 482722 630954
rect 482846 630854 482946 630954
rect 483070 630854 483170 630954
rect 482174 630630 482274 630730
rect 482398 630630 482498 630730
rect 482622 630630 482722 630730
rect 482846 630630 482946 630730
rect 483070 630630 483170 630730
rect 482174 630406 482274 630506
rect 482398 630406 482498 630506
rect 482622 630406 482722 630506
rect 482846 630406 482946 630506
rect 483070 630406 483170 630506
rect 482174 630182 482274 630282
rect 482398 630182 482498 630282
rect 482622 630182 482722 630282
rect 482846 630182 482946 630282
rect 483070 630182 483170 630282
rect 476352 630082 476404 630134
rect 476456 630082 476508 630134
rect 476560 630082 476612 630134
rect 476664 630082 476716 630134
rect 476768 630082 476820 630134
rect 476872 630082 476924 630134
rect 476352 629978 476404 630030
rect 476456 629978 476508 630030
rect 476560 629978 476612 630030
rect 476664 629978 476716 630030
rect 476768 629978 476820 630030
rect 476872 629978 476924 630030
rect 469218 629090 469358 629210
rect 454338 628930 454418 629010
rect 455258 628930 455338 629010
rect 456178 628930 456258 629010
rect 457098 628930 457178 629010
rect 458018 628930 458098 629010
rect 452848 628790 453248 628890
rect 459838 628930 459918 629010
rect 460758 628930 460838 629010
rect 461678 628930 461758 629010
rect 462598 628930 462678 629010
rect 463518 628930 463598 629010
rect 458758 628790 459158 628890
rect 465338 628930 465418 629010
rect 466258 628930 466338 629010
rect 467178 628930 467258 629010
rect 468098 628930 468178 629010
rect 469018 628930 469098 629010
rect 464258 628790 464658 628890
rect 470214 628788 470614 628888
rect 438920 627556 439020 627656
rect 439144 627556 439244 627656
rect 439368 627556 439468 627656
rect 439592 627556 439692 627656
rect 439816 627556 439916 627656
rect 440040 627556 440140 627656
rect 440264 627556 440364 627656
rect 440488 627556 440588 627656
rect 440712 627556 440812 627656
rect 440936 627556 441036 627656
rect 441160 627556 441260 627656
rect 441384 627556 441484 627656
rect 441608 627556 441708 627656
rect 441832 627556 441932 627656
rect 442056 627556 442156 627656
rect 442280 627556 442380 627656
rect 442504 627556 442604 627656
rect 442728 627556 442828 627656
rect 442952 627556 443052 627656
rect 443176 627556 443276 627656
rect 443400 627556 443500 627656
rect 443624 627556 443724 627656
rect 443848 627556 443948 627656
rect 444072 627556 444172 627656
rect 444296 627556 444396 627656
rect 444520 627556 444620 627656
rect 444744 627556 444844 627656
rect 444968 627556 445068 627656
rect 445192 627556 445292 627656
rect 445416 627556 445516 627656
rect 438920 627332 439020 627432
rect 439144 627332 439244 627432
rect 439368 627332 439468 627432
rect 439592 627332 439692 627432
rect 439816 627332 439916 627432
rect 440040 627332 440140 627432
rect 440264 627332 440364 627432
rect 440488 627332 440588 627432
rect 440712 627332 440812 627432
rect 440936 627332 441036 627432
rect 441160 627332 441260 627432
rect 441384 627332 441484 627432
rect 441608 627332 441708 627432
rect 441832 627332 441932 627432
rect 442056 627332 442156 627432
rect 442280 627332 442380 627432
rect 442504 627332 442604 627432
rect 442728 627332 442828 627432
rect 442952 627332 443052 627432
rect 443176 627332 443276 627432
rect 443400 627332 443500 627432
rect 443624 627332 443724 627432
rect 443848 627332 443948 627432
rect 444072 627332 444172 627432
rect 444296 627332 444396 627432
rect 444520 627332 444620 627432
rect 444744 627332 444844 627432
rect 444968 627332 445068 627432
rect 445192 627332 445292 627432
rect 445416 627332 445516 627432
rect 438920 627108 439020 627208
rect 439144 627108 439244 627208
rect 439368 627108 439468 627208
rect 439592 627108 439692 627208
rect 439816 627108 439916 627208
rect 440040 627108 440140 627208
rect 440264 627108 440364 627208
rect 440488 627108 440588 627208
rect 440712 627108 440812 627208
rect 440936 627108 441036 627208
rect 441160 627108 441260 627208
rect 441384 627108 441484 627208
rect 441608 627108 441708 627208
rect 441832 627108 441932 627208
rect 442056 627108 442156 627208
rect 442280 627108 442380 627208
rect 442504 627108 442604 627208
rect 442728 627108 442828 627208
rect 442952 627108 443052 627208
rect 443176 627108 443276 627208
rect 443400 627108 443500 627208
rect 443624 627108 443724 627208
rect 443848 627108 443948 627208
rect 444072 627108 444172 627208
rect 444296 627108 444396 627208
rect 444520 627108 444620 627208
rect 444744 627108 444844 627208
rect 444968 627108 445068 627208
rect 445192 627108 445292 627208
rect 445416 627108 445516 627208
rect 438920 626884 439020 626984
rect 439144 626884 439244 626984
rect 439368 626884 439468 626984
rect 439592 626884 439692 626984
rect 439816 626884 439916 626984
rect 440040 626884 440140 626984
rect 440264 626884 440364 626984
rect 440488 626884 440588 626984
rect 440712 626884 440812 626984
rect 440936 626884 441036 626984
rect 441160 626884 441260 626984
rect 441384 626884 441484 626984
rect 441608 626884 441708 626984
rect 441832 626884 441932 626984
rect 442056 626884 442156 626984
rect 442280 626884 442380 626984
rect 442504 626884 442604 626984
rect 442728 626884 442828 626984
rect 442952 626884 443052 626984
rect 443176 626884 443276 626984
rect 443400 626884 443500 626984
rect 443624 626884 443724 626984
rect 443848 626884 443948 626984
rect 444072 626884 444172 626984
rect 444296 626884 444396 626984
rect 444520 626884 444620 626984
rect 444744 626884 444844 626984
rect 444968 626884 445068 626984
rect 445192 626884 445292 626984
rect 445416 626884 445516 626984
rect 438920 626660 439020 626760
rect 439144 626660 439244 626760
rect 439368 626660 439468 626760
rect 439592 626660 439692 626760
rect 439816 626660 439916 626760
rect 440040 626660 440140 626760
rect 440264 626660 440364 626760
rect 440488 626660 440588 626760
rect 440712 626660 440812 626760
rect 440936 626660 441036 626760
rect 441160 626660 441260 626760
rect 441384 626660 441484 626760
rect 441608 626660 441708 626760
rect 441832 626660 441932 626760
rect 442056 626660 442156 626760
rect 442280 626660 442380 626760
rect 442504 626660 442604 626760
rect 442728 626660 442828 626760
rect 442952 626660 443052 626760
rect 443176 626660 443276 626760
rect 443400 626660 443500 626760
rect 443624 626660 443724 626760
rect 443848 626660 443948 626760
rect 444072 626660 444172 626760
rect 444296 626660 444396 626760
rect 444520 626660 444620 626760
rect 444744 626660 444844 626760
rect 444968 626660 445068 626760
rect 445192 626660 445292 626760
rect 445416 626660 445516 626760
rect 449390 627556 449490 627656
rect 449614 627556 449714 627656
rect 449838 627556 449938 627656
rect 450062 627556 450162 627656
rect 450286 627556 450386 627656
rect 450510 627556 450610 627656
rect 450734 627556 450834 627656
rect 450958 627556 451058 627656
rect 451182 627556 451282 627656
rect 451406 627556 451506 627656
rect 451630 627556 451730 627656
rect 451854 627556 451954 627656
rect 452078 627556 452178 627656
rect 452302 627556 452402 627656
rect 452526 627556 452626 627656
rect 452750 627556 452850 627656
rect 452974 627556 453074 627656
rect 453198 627556 453298 627656
rect 453422 627556 453522 627656
rect 453646 627556 453746 627656
rect 453870 627556 453970 627656
rect 454094 627556 454194 627656
rect 454318 627556 454418 627656
rect 454542 627556 454642 627656
rect 454766 627556 454866 627656
rect 454990 627556 455090 627656
rect 455214 627556 455314 627656
rect 455438 627556 455538 627656
rect 455662 627556 455762 627656
rect 455886 627556 455986 627656
rect 449390 627332 449490 627432
rect 449614 627332 449714 627432
rect 449838 627332 449938 627432
rect 450062 627332 450162 627432
rect 450286 627332 450386 627432
rect 450510 627332 450610 627432
rect 450734 627332 450834 627432
rect 450958 627332 451058 627432
rect 451182 627332 451282 627432
rect 451406 627332 451506 627432
rect 451630 627332 451730 627432
rect 451854 627332 451954 627432
rect 452078 627332 452178 627432
rect 452302 627332 452402 627432
rect 452526 627332 452626 627432
rect 452750 627332 452850 627432
rect 452974 627332 453074 627432
rect 453198 627332 453298 627432
rect 453422 627332 453522 627432
rect 453646 627332 453746 627432
rect 453870 627332 453970 627432
rect 454094 627332 454194 627432
rect 454318 627332 454418 627432
rect 454542 627332 454642 627432
rect 454766 627332 454866 627432
rect 454990 627332 455090 627432
rect 455214 627332 455314 627432
rect 455438 627332 455538 627432
rect 455662 627332 455762 627432
rect 455886 627332 455986 627432
rect 449390 627108 449490 627208
rect 449614 627108 449714 627208
rect 449838 627108 449938 627208
rect 450062 627108 450162 627208
rect 450286 627108 450386 627208
rect 450510 627108 450610 627208
rect 450734 627108 450834 627208
rect 450958 627108 451058 627208
rect 451182 627108 451282 627208
rect 451406 627108 451506 627208
rect 451630 627108 451730 627208
rect 451854 627108 451954 627208
rect 452078 627108 452178 627208
rect 452302 627108 452402 627208
rect 452526 627108 452626 627208
rect 452750 627108 452850 627208
rect 452974 627108 453074 627208
rect 453198 627108 453298 627208
rect 453422 627108 453522 627208
rect 453646 627108 453746 627208
rect 453870 627108 453970 627208
rect 454094 627108 454194 627208
rect 454318 627108 454418 627208
rect 454542 627108 454642 627208
rect 454766 627108 454866 627208
rect 454990 627108 455090 627208
rect 455214 627108 455314 627208
rect 455438 627108 455538 627208
rect 455662 627108 455762 627208
rect 455886 627108 455986 627208
rect 449390 626884 449490 626984
rect 449614 626884 449714 626984
rect 449838 626884 449938 626984
rect 450062 626884 450162 626984
rect 450286 626884 450386 626984
rect 450510 626884 450610 626984
rect 450734 626884 450834 626984
rect 450958 626884 451058 626984
rect 451182 626884 451282 626984
rect 451406 626884 451506 626984
rect 451630 626884 451730 626984
rect 451854 626884 451954 626984
rect 452078 626884 452178 626984
rect 452302 626884 452402 626984
rect 452526 626884 452626 626984
rect 452750 626884 452850 626984
rect 452974 626884 453074 626984
rect 453198 626884 453298 626984
rect 453422 626884 453522 626984
rect 453646 626884 453746 626984
rect 453870 626884 453970 626984
rect 454094 626884 454194 626984
rect 454318 626884 454418 626984
rect 454542 626884 454642 626984
rect 454766 626884 454866 626984
rect 454990 626884 455090 626984
rect 455214 626884 455314 626984
rect 455438 626884 455538 626984
rect 455662 626884 455762 626984
rect 455886 626884 455986 626984
rect 449390 626660 449490 626760
rect 449614 626660 449714 626760
rect 449838 626660 449938 626760
rect 450062 626660 450162 626760
rect 450286 626660 450386 626760
rect 450510 626660 450610 626760
rect 450734 626660 450834 626760
rect 450958 626660 451058 626760
rect 451182 626660 451282 626760
rect 451406 626660 451506 626760
rect 451630 626660 451730 626760
rect 451854 626660 451954 626760
rect 452078 626660 452178 626760
rect 452302 626660 452402 626760
rect 452526 626660 452626 626760
rect 452750 626660 452850 626760
rect 452974 626660 453074 626760
rect 453198 626660 453298 626760
rect 453422 626660 453522 626760
rect 453646 626660 453746 626760
rect 453870 626660 453970 626760
rect 454094 626660 454194 626760
rect 454318 626660 454418 626760
rect 454542 626660 454642 626760
rect 454766 626660 454866 626760
rect 454990 626660 455090 626760
rect 455214 626660 455314 626760
rect 455438 626660 455538 626760
rect 455662 626660 455762 626760
rect 455886 626660 455986 626760
rect 475660 627576 475760 627676
rect 475884 627576 475984 627676
rect 476108 627576 476208 627676
rect 476332 627576 476432 627676
rect 476556 627576 476656 627676
rect 476780 627576 476880 627676
rect 477004 627576 477104 627676
rect 477228 627576 477328 627676
rect 477452 627576 477552 627676
rect 477676 627576 477776 627676
rect 477900 627576 478000 627676
rect 478124 627576 478224 627676
rect 478348 627576 478448 627676
rect 478572 627576 478672 627676
rect 478796 627576 478896 627676
rect 479020 627576 479120 627676
rect 479244 627576 479344 627676
rect 479468 627576 479568 627676
rect 479692 627576 479792 627676
rect 479916 627576 480016 627676
rect 480140 627576 480240 627676
rect 480364 627576 480464 627676
rect 480588 627576 480688 627676
rect 480812 627576 480912 627676
rect 481036 627576 481136 627676
rect 481260 627576 481360 627676
rect 481484 627576 481584 627676
rect 481708 627576 481808 627676
rect 481932 627576 482032 627676
rect 482156 627576 482256 627676
rect 475660 627352 475760 627452
rect 475884 627352 475984 627452
rect 476108 627352 476208 627452
rect 476332 627352 476432 627452
rect 476556 627352 476656 627452
rect 476780 627352 476880 627452
rect 477004 627352 477104 627452
rect 477228 627352 477328 627452
rect 477452 627352 477552 627452
rect 477676 627352 477776 627452
rect 477900 627352 478000 627452
rect 478124 627352 478224 627452
rect 478348 627352 478448 627452
rect 478572 627352 478672 627452
rect 478796 627352 478896 627452
rect 479020 627352 479120 627452
rect 479244 627352 479344 627452
rect 479468 627352 479568 627452
rect 479692 627352 479792 627452
rect 479916 627352 480016 627452
rect 480140 627352 480240 627452
rect 480364 627352 480464 627452
rect 480588 627352 480688 627452
rect 480812 627352 480912 627452
rect 481036 627352 481136 627452
rect 481260 627352 481360 627452
rect 481484 627352 481584 627452
rect 481708 627352 481808 627452
rect 481932 627352 482032 627452
rect 482156 627352 482256 627452
rect 475660 627128 475760 627228
rect 475884 627128 475984 627228
rect 476108 627128 476208 627228
rect 476332 627128 476432 627228
rect 476556 627128 476656 627228
rect 476780 627128 476880 627228
rect 477004 627128 477104 627228
rect 477228 627128 477328 627228
rect 477452 627128 477552 627228
rect 477676 627128 477776 627228
rect 477900 627128 478000 627228
rect 478124 627128 478224 627228
rect 478348 627128 478448 627228
rect 478572 627128 478672 627228
rect 478796 627128 478896 627228
rect 479020 627128 479120 627228
rect 479244 627128 479344 627228
rect 479468 627128 479568 627228
rect 479692 627128 479792 627228
rect 479916 627128 480016 627228
rect 480140 627128 480240 627228
rect 480364 627128 480464 627228
rect 480588 627128 480688 627228
rect 480812 627128 480912 627228
rect 481036 627128 481136 627228
rect 481260 627128 481360 627228
rect 481484 627128 481584 627228
rect 481708 627128 481808 627228
rect 481932 627128 482032 627228
rect 482156 627128 482256 627228
rect 475660 626904 475760 627004
rect 475884 626904 475984 627004
rect 476108 626904 476208 627004
rect 476332 626904 476432 627004
rect 476556 626904 476656 627004
rect 476780 626904 476880 627004
rect 477004 626904 477104 627004
rect 477228 626904 477328 627004
rect 477452 626904 477552 627004
rect 477676 626904 477776 627004
rect 477900 626904 478000 627004
rect 478124 626904 478224 627004
rect 478348 626904 478448 627004
rect 478572 626904 478672 627004
rect 478796 626904 478896 627004
rect 479020 626904 479120 627004
rect 479244 626904 479344 627004
rect 479468 626904 479568 627004
rect 479692 626904 479792 627004
rect 479916 626904 480016 627004
rect 480140 626904 480240 627004
rect 480364 626904 480464 627004
rect 480588 626904 480688 627004
rect 480812 626904 480912 627004
rect 481036 626904 481136 627004
rect 481260 626904 481360 627004
rect 481484 626904 481584 627004
rect 481708 626904 481808 627004
rect 481932 626904 482032 627004
rect 482156 626904 482256 627004
rect 475660 626680 475760 626780
rect 475884 626680 475984 626780
rect 476108 626680 476208 626780
rect 476332 626680 476432 626780
rect 476556 626680 476656 626780
rect 476780 626680 476880 626780
rect 477004 626680 477104 626780
rect 477228 626680 477328 626780
rect 477452 626680 477552 626780
rect 477676 626680 477776 626780
rect 477900 626680 478000 626780
rect 478124 626680 478224 626780
rect 478348 626680 478448 626780
rect 478572 626680 478672 626780
rect 478796 626680 478896 626780
rect 479020 626680 479120 626780
rect 479244 626680 479344 626780
rect 479468 626680 479568 626780
rect 479692 626680 479792 626780
rect 479916 626680 480016 626780
rect 480140 626680 480240 626780
rect 480364 626680 480464 626780
rect 480588 626680 480688 626780
rect 480812 626680 480912 626780
rect 481036 626680 481136 626780
rect 481260 626680 481360 626780
rect 481484 626680 481584 626780
rect 481708 626680 481808 626780
rect 481932 626680 482032 626780
rect 482156 626680 482256 626780
<< metal2 >>
rect 438880 654876 445540 654906
rect 438880 654776 438920 654876
rect 439020 654776 439144 654876
rect 439244 654776 439368 654876
rect 439468 654776 439592 654876
rect 439692 654776 439816 654876
rect 439916 654776 440040 654876
rect 440140 654776 440264 654876
rect 440364 654776 440488 654876
rect 440588 654776 440712 654876
rect 440812 654776 440936 654876
rect 441036 654776 441160 654876
rect 441260 654776 441384 654876
rect 441484 654776 441608 654876
rect 441708 654776 441832 654876
rect 441932 654776 442056 654876
rect 442156 654776 442280 654876
rect 442380 654776 442504 654876
rect 442604 654776 442728 654876
rect 442828 654776 442952 654876
rect 443052 654776 443176 654876
rect 443276 654776 443400 654876
rect 443500 654776 443624 654876
rect 443724 654776 443848 654876
rect 443948 654776 444072 654876
rect 444172 654776 444296 654876
rect 444396 654776 444520 654876
rect 444620 654776 444744 654876
rect 444844 654776 444968 654876
rect 445068 654776 445192 654876
rect 445292 654776 445416 654876
rect 445516 654776 445540 654876
rect 438880 654652 445540 654776
rect 438880 654552 438920 654652
rect 439020 654552 439144 654652
rect 439244 654552 439368 654652
rect 439468 654552 439592 654652
rect 439692 654552 439816 654652
rect 439916 654552 440040 654652
rect 440140 654552 440264 654652
rect 440364 654552 440488 654652
rect 440588 654552 440712 654652
rect 440812 654552 440936 654652
rect 441036 654552 441160 654652
rect 441260 654552 441384 654652
rect 441484 654552 441608 654652
rect 441708 654552 441832 654652
rect 441932 654552 442056 654652
rect 442156 654552 442280 654652
rect 442380 654552 442504 654652
rect 442604 654552 442728 654652
rect 442828 654552 442952 654652
rect 443052 654552 443176 654652
rect 443276 654552 443400 654652
rect 443500 654552 443624 654652
rect 443724 654552 443848 654652
rect 443948 654552 444072 654652
rect 444172 654552 444296 654652
rect 444396 654552 444520 654652
rect 444620 654552 444744 654652
rect 444844 654552 444968 654652
rect 445068 654552 445192 654652
rect 445292 654552 445416 654652
rect 445516 654552 445540 654652
rect 438880 654428 445540 654552
rect 438880 654328 438920 654428
rect 439020 654328 439144 654428
rect 439244 654328 439368 654428
rect 439468 654328 439592 654428
rect 439692 654328 439816 654428
rect 439916 654328 440040 654428
rect 440140 654328 440264 654428
rect 440364 654328 440488 654428
rect 440588 654328 440712 654428
rect 440812 654328 440936 654428
rect 441036 654328 441160 654428
rect 441260 654328 441384 654428
rect 441484 654328 441608 654428
rect 441708 654328 441832 654428
rect 441932 654328 442056 654428
rect 442156 654328 442280 654428
rect 442380 654328 442504 654428
rect 442604 654328 442728 654428
rect 442828 654328 442952 654428
rect 443052 654328 443176 654428
rect 443276 654328 443400 654428
rect 443500 654328 443624 654428
rect 443724 654328 443848 654428
rect 443948 654328 444072 654428
rect 444172 654328 444296 654428
rect 444396 654328 444520 654428
rect 444620 654328 444744 654428
rect 444844 654328 444968 654428
rect 445068 654328 445192 654428
rect 445292 654328 445416 654428
rect 445516 654328 445540 654428
rect 438880 654204 445540 654328
rect 438880 654104 438920 654204
rect 439020 654104 439144 654204
rect 439244 654104 439368 654204
rect 439468 654104 439592 654204
rect 439692 654104 439816 654204
rect 439916 654104 440040 654204
rect 440140 654104 440264 654204
rect 440364 654104 440488 654204
rect 440588 654104 440712 654204
rect 440812 654104 440936 654204
rect 441036 654104 441160 654204
rect 441260 654104 441384 654204
rect 441484 654104 441608 654204
rect 441708 654104 441832 654204
rect 441932 654104 442056 654204
rect 442156 654104 442280 654204
rect 442380 654104 442504 654204
rect 442604 654104 442728 654204
rect 442828 654104 442952 654204
rect 443052 654104 443176 654204
rect 443276 654104 443400 654204
rect 443500 654104 443624 654204
rect 443724 654104 443848 654204
rect 443948 654104 444072 654204
rect 444172 654104 444296 654204
rect 444396 654104 444520 654204
rect 444620 654104 444744 654204
rect 444844 654104 444968 654204
rect 445068 654104 445192 654204
rect 445292 654104 445416 654204
rect 445516 654104 445540 654204
rect 438880 653980 445540 654104
rect 438880 653880 438920 653980
rect 439020 653880 439144 653980
rect 439244 653880 439368 653980
rect 439468 653880 439592 653980
rect 439692 653880 439816 653980
rect 439916 653880 440040 653980
rect 440140 653880 440264 653980
rect 440364 653880 440488 653980
rect 440588 653880 440712 653980
rect 440812 653880 440936 653980
rect 441036 653880 441160 653980
rect 441260 653880 441384 653980
rect 441484 653880 441608 653980
rect 441708 653880 441832 653980
rect 441932 653880 442056 653980
rect 442156 653880 442280 653980
rect 442380 653880 442504 653980
rect 442604 653880 442728 653980
rect 442828 653880 442952 653980
rect 443052 653880 443176 653980
rect 443276 653880 443400 653980
rect 443500 653880 443624 653980
rect 443724 653880 443848 653980
rect 443948 653880 444072 653980
rect 444172 653880 444296 653980
rect 444396 653880 444520 653980
rect 444620 653880 444744 653980
rect 444844 653880 444968 653980
rect 445068 653880 445192 653980
rect 445292 653880 445416 653980
rect 445516 653880 445540 653980
rect 438880 653846 445540 653880
rect 449350 654876 456010 654906
rect 449350 654776 449390 654876
rect 449490 654776 449614 654876
rect 449714 654776 449838 654876
rect 449938 654776 450062 654876
rect 450162 654776 450286 654876
rect 450386 654776 450510 654876
rect 450610 654776 450734 654876
rect 450834 654776 450958 654876
rect 451058 654776 451182 654876
rect 451282 654776 451406 654876
rect 451506 654776 451630 654876
rect 451730 654776 451854 654876
rect 451954 654776 452078 654876
rect 452178 654776 452302 654876
rect 452402 654776 452526 654876
rect 452626 654776 452750 654876
rect 452850 654776 452974 654876
rect 453074 654776 453198 654876
rect 453298 654776 453422 654876
rect 453522 654776 453646 654876
rect 453746 654776 453870 654876
rect 453970 654776 454094 654876
rect 454194 654776 454318 654876
rect 454418 654776 454542 654876
rect 454642 654776 454766 654876
rect 454866 654776 454990 654876
rect 455090 654776 455214 654876
rect 455314 654776 455438 654876
rect 455538 654776 455662 654876
rect 455762 654776 455886 654876
rect 455986 654776 456010 654876
rect 449350 654652 456010 654776
rect 449350 654552 449390 654652
rect 449490 654552 449614 654652
rect 449714 654552 449838 654652
rect 449938 654552 450062 654652
rect 450162 654552 450286 654652
rect 450386 654552 450510 654652
rect 450610 654552 450734 654652
rect 450834 654552 450958 654652
rect 451058 654552 451182 654652
rect 451282 654552 451406 654652
rect 451506 654552 451630 654652
rect 451730 654552 451854 654652
rect 451954 654552 452078 654652
rect 452178 654552 452302 654652
rect 452402 654552 452526 654652
rect 452626 654552 452750 654652
rect 452850 654552 452974 654652
rect 453074 654552 453198 654652
rect 453298 654552 453422 654652
rect 453522 654552 453646 654652
rect 453746 654552 453870 654652
rect 453970 654552 454094 654652
rect 454194 654552 454318 654652
rect 454418 654552 454542 654652
rect 454642 654552 454766 654652
rect 454866 654552 454990 654652
rect 455090 654552 455214 654652
rect 455314 654552 455438 654652
rect 455538 654552 455662 654652
rect 455762 654552 455886 654652
rect 455986 654552 456010 654652
rect 449350 654428 456010 654552
rect 449350 654328 449390 654428
rect 449490 654328 449614 654428
rect 449714 654328 449838 654428
rect 449938 654328 450062 654428
rect 450162 654328 450286 654428
rect 450386 654328 450510 654428
rect 450610 654328 450734 654428
rect 450834 654328 450958 654428
rect 451058 654328 451182 654428
rect 451282 654328 451406 654428
rect 451506 654328 451630 654428
rect 451730 654328 451854 654428
rect 451954 654328 452078 654428
rect 452178 654328 452302 654428
rect 452402 654328 452526 654428
rect 452626 654328 452750 654428
rect 452850 654328 452974 654428
rect 453074 654328 453198 654428
rect 453298 654328 453422 654428
rect 453522 654328 453646 654428
rect 453746 654328 453870 654428
rect 453970 654328 454094 654428
rect 454194 654328 454318 654428
rect 454418 654328 454542 654428
rect 454642 654328 454766 654428
rect 454866 654328 454990 654428
rect 455090 654328 455214 654428
rect 455314 654328 455438 654428
rect 455538 654328 455662 654428
rect 455762 654328 455886 654428
rect 455986 654328 456010 654428
rect 449350 654204 456010 654328
rect 449350 654104 449390 654204
rect 449490 654104 449614 654204
rect 449714 654104 449838 654204
rect 449938 654104 450062 654204
rect 450162 654104 450286 654204
rect 450386 654104 450510 654204
rect 450610 654104 450734 654204
rect 450834 654104 450958 654204
rect 451058 654104 451182 654204
rect 451282 654104 451406 654204
rect 451506 654104 451630 654204
rect 451730 654104 451854 654204
rect 451954 654104 452078 654204
rect 452178 654104 452302 654204
rect 452402 654104 452526 654204
rect 452626 654104 452750 654204
rect 452850 654104 452974 654204
rect 453074 654104 453198 654204
rect 453298 654104 453422 654204
rect 453522 654104 453646 654204
rect 453746 654104 453870 654204
rect 453970 654104 454094 654204
rect 454194 654104 454318 654204
rect 454418 654104 454542 654204
rect 454642 654104 454766 654204
rect 454866 654104 454990 654204
rect 455090 654104 455214 654204
rect 455314 654104 455438 654204
rect 455538 654104 455662 654204
rect 455762 654104 455886 654204
rect 455986 654104 456010 654204
rect 449350 653980 456010 654104
rect 449350 653880 449390 653980
rect 449490 653880 449614 653980
rect 449714 653880 449838 653980
rect 449938 653880 450062 653980
rect 450162 653880 450286 653980
rect 450386 653880 450510 653980
rect 450610 653880 450734 653980
rect 450834 653880 450958 653980
rect 451058 653880 451182 653980
rect 451282 653880 451406 653980
rect 451506 653880 451630 653980
rect 451730 653880 451854 653980
rect 451954 653880 452078 653980
rect 452178 653880 452302 653980
rect 452402 653880 452526 653980
rect 452626 653880 452750 653980
rect 452850 653880 452974 653980
rect 453074 653880 453198 653980
rect 453298 653880 453422 653980
rect 453522 653880 453646 653980
rect 453746 653880 453870 653980
rect 453970 653880 454094 653980
rect 454194 653880 454318 653980
rect 454418 653880 454542 653980
rect 454642 653880 454766 653980
rect 454866 653880 454990 653980
rect 455090 653880 455214 653980
rect 455314 653880 455438 653980
rect 455538 653880 455662 653980
rect 455762 653880 455886 653980
rect 455986 653880 456010 653980
rect 449350 653846 456010 653880
rect 475620 654896 482280 654926
rect 475620 654796 475660 654896
rect 475760 654796 475884 654896
rect 475984 654796 476108 654896
rect 476208 654796 476332 654896
rect 476432 654796 476556 654896
rect 476656 654796 476780 654896
rect 476880 654796 477004 654896
rect 477104 654796 477228 654896
rect 477328 654796 477452 654896
rect 477552 654796 477676 654896
rect 477776 654796 477900 654896
rect 478000 654796 478124 654896
rect 478224 654796 478348 654896
rect 478448 654796 478572 654896
rect 478672 654796 478796 654896
rect 478896 654796 479020 654896
rect 479120 654796 479244 654896
rect 479344 654796 479468 654896
rect 479568 654796 479692 654896
rect 479792 654796 479916 654896
rect 480016 654796 480140 654896
rect 480240 654796 480364 654896
rect 480464 654796 480588 654896
rect 480688 654796 480812 654896
rect 480912 654796 481036 654896
rect 481136 654796 481260 654896
rect 481360 654796 481484 654896
rect 481584 654796 481708 654896
rect 481808 654796 481932 654896
rect 482032 654796 482156 654896
rect 482256 654796 482280 654896
rect 475620 654672 482280 654796
rect 475620 654572 475660 654672
rect 475760 654572 475884 654672
rect 475984 654572 476108 654672
rect 476208 654572 476332 654672
rect 476432 654572 476556 654672
rect 476656 654572 476780 654672
rect 476880 654572 477004 654672
rect 477104 654572 477228 654672
rect 477328 654572 477452 654672
rect 477552 654572 477676 654672
rect 477776 654572 477900 654672
rect 478000 654572 478124 654672
rect 478224 654572 478348 654672
rect 478448 654572 478572 654672
rect 478672 654572 478796 654672
rect 478896 654572 479020 654672
rect 479120 654572 479244 654672
rect 479344 654572 479468 654672
rect 479568 654572 479692 654672
rect 479792 654572 479916 654672
rect 480016 654572 480140 654672
rect 480240 654572 480364 654672
rect 480464 654572 480588 654672
rect 480688 654572 480812 654672
rect 480912 654572 481036 654672
rect 481136 654572 481260 654672
rect 481360 654572 481484 654672
rect 481584 654572 481708 654672
rect 481808 654572 481932 654672
rect 482032 654572 482156 654672
rect 482256 654572 482280 654672
rect 475620 654448 482280 654572
rect 475620 654348 475660 654448
rect 475760 654348 475884 654448
rect 475984 654348 476108 654448
rect 476208 654348 476332 654448
rect 476432 654348 476556 654448
rect 476656 654348 476780 654448
rect 476880 654348 477004 654448
rect 477104 654348 477228 654448
rect 477328 654348 477452 654448
rect 477552 654348 477676 654448
rect 477776 654348 477900 654448
rect 478000 654348 478124 654448
rect 478224 654348 478348 654448
rect 478448 654348 478572 654448
rect 478672 654348 478796 654448
rect 478896 654348 479020 654448
rect 479120 654348 479244 654448
rect 479344 654348 479468 654448
rect 479568 654348 479692 654448
rect 479792 654348 479916 654448
rect 480016 654348 480140 654448
rect 480240 654348 480364 654448
rect 480464 654348 480588 654448
rect 480688 654348 480812 654448
rect 480912 654348 481036 654448
rect 481136 654348 481260 654448
rect 481360 654348 481484 654448
rect 481584 654348 481708 654448
rect 481808 654348 481932 654448
rect 482032 654348 482156 654448
rect 482256 654348 482280 654448
rect 475620 654224 482280 654348
rect 475620 654124 475660 654224
rect 475760 654124 475884 654224
rect 475984 654124 476108 654224
rect 476208 654124 476332 654224
rect 476432 654124 476556 654224
rect 476656 654124 476780 654224
rect 476880 654124 477004 654224
rect 477104 654124 477228 654224
rect 477328 654124 477452 654224
rect 477552 654124 477676 654224
rect 477776 654124 477900 654224
rect 478000 654124 478124 654224
rect 478224 654124 478348 654224
rect 478448 654124 478572 654224
rect 478672 654124 478796 654224
rect 478896 654124 479020 654224
rect 479120 654124 479244 654224
rect 479344 654124 479468 654224
rect 479568 654124 479692 654224
rect 479792 654124 479916 654224
rect 480016 654124 480140 654224
rect 480240 654124 480364 654224
rect 480464 654124 480588 654224
rect 480688 654124 480812 654224
rect 480912 654124 481036 654224
rect 481136 654124 481260 654224
rect 481360 654124 481484 654224
rect 481584 654124 481708 654224
rect 481808 654124 481932 654224
rect 482032 654124 482156 654224
rect 482256 654124 482280 654224
rect 475620 654000 482280 654124
rect 475620 653900 475660 654000
rect 475760 653900 475884 654000
rect 475984 653900 476108 654000
rect 476208 653900 476332 654000
rect 476432 653900 476556 654000
rect 476656 653900 476780 654000
rect 476880 653900 477004 654000
rect 477104 653900 477228 654000
rect 477328 653900 477452 654000
rect 477552 653900 477676 654000
rect 477776 653900 477900 654000
rect 478000 653900 478124 654000
rect 478224 653900 478348 654000
rect 478448 653900 478572 654000
rect 478672 653900 478796 654000
rect 478896 653900 479020 654000
rect 479120 653900 479244 654000
rect 479344 653900 479468 654000
rect 479568 653900 479692 654000
rect 479792 653900 479916 654000
rect 480016 653900 480140 654000
rect 480240 653900 480364 654000
rect 480464 653900 480588 654000
rect 480688 653900 480812 654000
rect 480912 653900 481036 654000
rect 481136 653900 481260 654000
rect 481360 653900 481484 654000
rect 481584 653900 481708 654000
rect 481808 653900 481932 654000
rect 482032 653900 482156 654000
rect 482256 653900 482280 654000
rect 475620 653866 482280 653900
rect 440687 652760 451961 652769
rect 440687 651922 440696 652760
rect 451952 651922 451961 652760
rect 440687 651913 451961 651922
rect 463962 651214 464532 651220
rect 463962 650656 463968 651214
rect 464526 650656 464532 651214
rect 457406 650414 457976 650420
rect 437864 650178 438924 650202
rect 437864 650078 437894 650178
rect 437994 650078 438118 650178
rect 438218 650078 438342 650178
rect 438442 650078 438566 650178
rect 438666 650078 438790 650178
rect 438890 650078 438924 650178
rect 437864 649954 438924 650078
rect 437864 649854 437894 649954
rect 437994 649854 438118 649954
rect 438218 649854 438342 649954
rect 438442 649854 438566 649954
rect 438666 649854 438790 649954
rect 438890 649854 438924 649954
rect 437864 649730 438924 649854
rect 437864 649630 437894 649730
rect 437994 649630 438118 649730
rect 438218 649630 438342 649730
rect 438442 649630 438566 649730
rect 438666 649630 438790 649730
rect 438890 649630 438924 649730
rect 437864 649506 438924 649630
rect 437864 649406 437894 649506
rect 437994 649406 438118 649506
rect 438218 649406 438342 649506
rect 438442 649406 438566 649506
rect 438666 649406 438790 649506
rect 438890 649406 438924 649506
rect 437864 649282 438924 649406
rect 437864 649182 437894 649282
rect 437994 649182 438118 649282
rect 438218 649182 438342 649282
rect 438442 649182 438566 649282
rect 438666 649182 438790 649282
rect 438890 649182 438924 649282
rect 457406 649856 457412 650414
rect 457970 649856 457976 650414
rect 457406 649676 457976 649856
rect 463132 650414 463702 650420
rect 463132 649856 463138 650414
rect 463696 649856 463702 650414
rect 457406 649256 457412 649676
rect 457970 649256 457976 649676
rect 457406 649250 457976 649256
rect 458224 649676 458794 649682
rect 458224 649256 458230 649676
rect 458788 649256 458794 649676
rect 437864 649058 438924 649182
rect 437864 648958 437894 649058
rect 437994 648958 438118 649058
rect 438218 648958 438342 649058
rect 438442 648958 438566 649058
rect 438666 648958 438790 649058
rect 438890 648958 438924 649058
rect 437864 648834 438924 648958
rect 437864 648734 437894 648834
rect 437994 648734 438118 648834
rect 438218 648734 438342 648834
rect 438442 648734 438566 648834
rect 438666 648734 438790 648834
rect 438890 648734 438924 648834
rect 437864 648610 438924 648734
rect 437864 648510 437894 648610
rect 437994 648510 438118 648610
rect 438218 648510 438342 648610
rect 438442 648510 438566 648610
rect 438666 648510 438790 648610
rect 438890 648510 438924 648610
rect 437864 648386 438924 648510
rect 458224 648952 458794 649256
rect 458224 648460 458230 648952
rect 458788 648460 458794 648952
rect 458224 648450 458794 648460
rect 462314 649614 462884 649620
rect 462314 649194 462320 649614
rect 462878 649194 462884 649614
rect 462314 648952 462884 649194
rect 463132 649614 463702 649856
rect 463962 649620 464532 650656
rect 465586 651214 466156 651220
rect 465586 650656 465592 651214
rect 466150 650656 466156 651214
rect 463132 649194 463138 649614
rect 463696 649194 463702 649614
rect 463132 649188 463702 649194
rect 463950 649614 464532 649620
rect 463950 649194 463956 649614
rect 464514 649206 464532 649614
rect 464768 649614 465338 649620
rect 464514 649194 464520 649206
rect 463950 649188 464520 649194
rect 464768 649194 464774 649614
rect 465332 649194 465338 649614
rect 462314 648394 462320 648952
rect 462878 648394 462884 648952
rect 462314 648388 462884 648394
rect 464768 648952 465338 649194
rect 465586 649614 466156 650656
rect 469676 651214 470246 651220
rect 469676 650656 469682 651214
rect 470240 650656 470246 651214
rect 465586 649194 465592 649614
rect 466150 649194 466156 649614
rect 465586 649188 466156 649194
rect 466404 650414 466974 650420
rect 466404 649856 466410 650414
rect 466968 649856 466974 650414
rect 466404 649614 466974 649856
rect 468858 650414 469428 650420
rect 468858 649856 468864 650414
rect 469422 649856 469428 650414
rect 466404 649194 466410 649614
rect 466968 649194 466974 649614
rect 466404 649188 466974 649194
rect 467222 649614 467792 649620
rect 467222 649194 467228 649614
rect 467786 649194 467792 649614
rect 464768 648394 464774 648952
rect 465332 648394 465338 648952
rect 464768 648388 465338 648394
rect 467222 648952 467792 649194
rect 467222 648394 467228 648952
rect 467786 648394 467792 648952
rect 467222 648388 467792 648394
rect 468040 649614 468610 649620
rect 468040 649194 468046 649614
rect 468604 649194 468610 649614
rect 437864 648286 437894 648386
rect 437994 648286 438118 648386
rect 438218 648286 438342 648386
rect 438442 648286 438566 648386
rect 438666 648286 438790 648386
rect 438890 648286 438924 648386
rect 437864 648162 438924 648286
rect 437864 648062 437894 648162
rect 437994 648062 438118 648162
rect 438218 648062 438342 648162
rect 438442 648062 438566 648162
rect 438666 648062 438790 648162
rect 438890 648062 438924 648162
rect 437864 647938 438924 648062
rect 437864 647838 437894 647938
rect 437994 647838 438118 647938
rect 438218 647838 438342 647938
rect 438442 647838 438566 647938
rect 438666 647838 438790 647938
rect 438890 647838 438924 647938
rect 437864 647714 438924 647838
rect 437864 647614 437894 647714
rect 437994 647614 438118 647714
rect 438218 647614 438342 647714
rect 438442 647614 438566 647714
rect 438666 647614 438790 647714
rect 438890 647614 438924 647714
rect 437864 647490 438924 647614
rect 437864 647390 437894 647490
rect 437994 647390 438118 647490
rect 438218 647390 438342 647490
rect 438442 647390 438566 647490
rect 438666 647390 438790 647490
rect 438890 647390 438924 647490
rect 437864 647266 438924 647390
rect 437864 647166 437894 647266
rect 437994 647166 438118 647266
rect 438218 647166 438342 647266
rect 438442 647166 438566 647266
rect 438666 647166 438790 647266
rect 438890 647166 438924 647266
rect 437864 647042 438924 647166
rect 437864 646942 437894 647042
rect 437994 646942 438118 647042
rect 438218 646942 438342 647042
rect 438442 646942 438566 647042
rect 438666 646942 438790 647042
rect 438890 646942 438924 647042
rect 437864 646818 438924 646942
rect 437864 646718 437894 646818
rect 437994 646718 438118 646818
rect 438218 646718 438342 646818
rect 438442 646718 438566 646818
rect 438666 646718 438790 646818
rect 438890 646718 438924 646818
rect 437864 646594 438924 646718
rect 437864 646494 437894 646594
rect 437994 646494 438118 646594
rect 438218 646494 438342 646594
rect 438442 646494 438566 646594
rect 438666 646494 438790 646594
rect 438890 646494 438924 646594
rect 437864 646370 438924 646494
rect 437864 646270 437894 646370
rect 437994 646270 438118 646370
rect 438218 646270 438342 646370
rect 438442 646270 438566 646370
rect 438666 646270 438790 646370
rect 438890 646270 438924 646370
rect 437864 646146 438924 646270
rect 468040 646758 468610 649194
rect 468858 649614 469428 649856
rect 468858 649194 468864 649614
rect 469422 649194 469428 649614
rect 468858 649188 469428 649194
rect 469676 649614 470246 650656
rect 472136 651214 472700 651220
rect 472694 650656 472700 651214
rect 472136 650650 472700 650656
rect 471312 650414 471882 650420
rect 471312 649856 471318 650414
rect 471876 649856 471882 650414
rect 469676 649194 469682 649614
rect 470240 649194 470246 649614
rect 469676 649188 470246 649194
rect 470494 649614 471064 649620
rect 470494 649194 470500 649614
rect 471058 649194 471064 649614
rect 470494 648952 471064 649194
rect 471312 649614 471882 649856
rect 471312 649194 471318 649614
rect 471876 649194 471882 649614
rect 471312 649188 471882 649194
rect 472130 649614 472700 650650
rect 473766 650414 474336 650420
rect 473766 649856 473772 650414
rect 474330 649856 474336 650414
rect 472130 649194 472136 649614
rect 472694 649194 472700 649614
rect 472130 649188 472700 649194
rect 472948 649614 473518 649620
rect 472948 649194 472954 649614
rect 473512 649194 473518 649614
rect 470494 648394 470500 648952
rect 471058 648394 471064 648952
rect 470494 648388 471064 648394
rect 472948 648952 473518 649194
rect 473766 649614 474336 649856
rect 473766 649194 473772 649614
rect 474330 649194 474336 649614
rect 473766 649188 474336 649194
rect 482144 650178 483204 650202
rect 482144 650078 482174 650178
rect 482274 650078 482398 650178
rect 482498 650078 482622 650178
rect 482722 650078 482846 650178
rect 482946 650078 483070 650178
rect 483170 650078 483204 650178
rect 482144 649954 483204 650078
rect 482144 649854 482174 649954
rect 482274 649854 482398 649954
rect 482498 649854 482622 649954
rect 482722 649854 482846 649954
rect 482946 649854 483070 649954
rect 483170 649854 483204 649954
rect 482144 649730 483204 649854
rect 482144 649630 482174 649730
rect 482274 649630 482398 649730
rect 482498 649630 482622 649730
rect 482722 649630 482846 649730
rect 482946 649630 483070 649730
rect 483170 649630 483204 649730
rect 482144 649506 483204 649630
rect 482144 649406 482174 649506
rect 482274 649406 482398 649506
rect 482498 649406 482622 649506
rect 482722 649406 482846 649506
rect 482946 649406 483070 649506
rect 483170 649406 483204 649506
rect 482144 649282 483204 649406
rect 472948 648394 472954 648952
rect 473512 648394 473518 648952
rect 472948 648388 473518 648394
rect 482144 649182 482174 649282
rect 482274 649182 482398 649282
rect 482498 649182 482622 649282
rect 482722 649182 482846 649282
rect 482946 649182 483070 649282
rect 483170 649182 483204 649282
rect 482144 649058 483204 649182
rect 482144 648958 482174 649058
rect 482274 648958 482398 649058
rect 482498 648958 482622 649058
rect 482722 648958 482846 649058
rect 482946 648958 483070 649058
rect 483170 648958 483204 649058
rect 482144 648834 483204 648958
rect 482144 648734 482174 648834
rect 482274 648734 482398 648834
rect 482498 648734 482622 648834
rect 482722 648734 482846 648834
rect 482946 648734 483070 648834
rect 483170 648734 483204 648834
rect 482144 648610 483204 648734
rect 482144 648510 482174 648610
rect 482274 648510 482398 648610
rect 482498 648510 482622 648610
rect 482722 648510 482846 648610
rect 482946 648510 483070 648610
rect 483170 648510 483204 648610
rect 482144 648386 483204 648510
rect 482144 648286 482174 648386
rect 482274 648286 482398 648386
rect 482498 648286 482622 648386
rect 482722 648286 482846 648386
rect 482946 648286 483070 648386
rect 483170 648286 483204 648386
rect 482144 648162 483204 648286
rect 482144 648062 482174 648162
rect 482274 648062 482398 648162
rect 482498 648062 482622 648162
rect 482722 648062 482846 648162
rect 482946 648062 483070 648162
rect 483170 648062 483204 648162
rect 482144 647938 483204 648062
rect 482144 647838 482174 647938
rect 482274 647838 482398 647938
rect 482498 647838 482622 647938
rect 482722 647838 482846 647938
rect 482946 647838 483070 647938
rect 483170 647838 483204 647938
rect 482144 647714 483204 647838
rect 482144 647614 482174 647714
rect 482274 647614 482398 647714
rect 482498 647614 482622 647714
rect 482722 647614 482846 647714
rect 482946 647614 483070 647714
rect 483170 647614 483204 647714
rect 482144 647490 483204 647614
rect 482144 647390 482174 647490
rect 482274 647390 482398 647490
rect 482498 647390 482622 647490
rect 482722 647390 482846 647490
rect 482946 647390 483070 647490
rect 483170 647390 483204 647490
rect 482144 647266 483204 647390
rect 482144 647166 482174 647266
rect 482274 647166 482398 647266
rect 482498 647166 482622 647266
rect 482722 647166 482846 647266
rect 482946 647166 483070 647266
rect 483170 647166 483204 647266
rect 482144 647042 483204 647166
rect 482144 646942 482174 647042
rect 482274 646942 482398 647042
rect 482498 646942 482622 647042
rect 482722 646942 482846 647042
rect 482946 646942 483070 647042
rect 483170 646942 483204 647042
rect 482144 646818 483204 646942
rect 468040 646188 474324 646758
rect 437864 646046 437894 646146
rect 437994 646046 438118 646146
rect 438218 646046 438342 646146
rect 438442 646046 438566 646146
rect 438666 646046 438790 646146
rect 438890 646046 438924 646146
rect 437864 645922 438924 646046
rect 437864 645822 437894 645922
rect 437994 645822 438118 645922
rect 438218 645822 438342 645922
rect 438442 645822 438566 645922
rect 438666 645822 438790 645922
rect 438890 645822 438924 645922
rect 437864 645698 438924 645822
rect 437864 645598 437894 645698
rect 437994 645598 438118 645698
rect 438218 645598 438342 645698
rect 438442 645598 438566 645698
rect 438666 645598 438790 645698
rect 438890 645598 438924 645698
rect 437864 645474 438924 645598
rect 437864 645374 437894 645474
rect 437994 645374 438118 645474
rect 438218 645374 438342 645474
rect 438442 645374 438566 645474
rect 438666 645374 438790 645474
rect 438890 645374 438924 645474
rect 437864 645250 438924 645374
rect 437864 645150 437894 645250
rect 437994 645150 438118 645250
rect 438218 645150 438342 645250
rect 438442 645150 438566 645250
rect 438666 645150 438790 645250
rect 438890 645150 438924 645250
rect 437864 645026 438924 645150
rect 437864 644926 437894 645026
rect 437994 644926 438118 645026
rect 438218 644926 438342 645026
rect 438442 644926 438566 645026
rect 438666 644926 438790 645026
rect 438890 644926 438924 645026
rect 437864 644802 438924 644926
rect 437864 644702 437894 644802
rect 437994 644702 438118 644802
rect 438218 644702 438342 644802
rect 438442 644702 438566 644802
rect 438666 644702 438790 644802
rect 438890 644702 438924 644802
rect 437864 644578 438924 644702
rect 437864 644478 437894 644578
rect 437994 644478 438118 644578
rect 438218 644478 438342 644578
rect 438442 644478 438566 644578
rect 438666 644478 438790 644578
rect 438890 644478 438924 644578
rect 437864 644354 438924 644478
rect 437864 644254 437894 644354
rect 437994 644254 438118 644354
rect 438218 644254 438342 644354
rect 438442 644254 438566 644354
rect 438666 644254 438790 644354
rect 438890 644254 438924 644354
rect 437864 644130 438924 644254
rect 437864 644030 437894 644130
rect 437994 644030 438118 644130
rect 438218 644030 438342 644130
rect 438442 644030 438566 644130
rect 438666 644030 438790 644130
rect 438890 644030 438924 644130
rect 437864 643906 438924 644030
rect 437864 643806 437894 643906
rect 437994 643806 438118 643906
rect 438218 643806 438342 643906
rect 438442 643806 438566 643906
rect 438666 643806 438790 643906
rect 438890 643806 438924 643906
rect 437864 643682 438924 643806
rect 437864 643582 437894 643682
rect 437994 643582 438118 643682
rect 438218 643582 438342 643682
rect 438442 643582 438566 643682
rect 438666 643582 438790 643682
rect 438890 643582 438924 643682
rect 437864 643542 438924 643582
rect 463132 644478 463702 644484
rect 463132 643920 463138 644478
rect 463696 643920 463702 644478
rect 462314 642878 462884 642884
rect 462314 642458 462320 642878
rect 462878 642458 462884 642878
rect 462314 642216 462884 642458
rect 463132 642878 463702 643920
rect 466404 644478 466974 644484
rect 466404 643920 466410 644478
rect 466968 643920 466974 644478
rect 463132 642458 463138 642878
rect 463696 642458 463702 642878
rect 463132 642452 463702 642458
rect 463950 643678 464520 643684
rect 463950 643120 463956 643678
rect 464514 643120 464520 643678
rect 463950 642878 464520 643120
rect 465586 643678 466156 643684
rect 465586 643120 465592 643678
rect 466150 643120 466156 643678
rect 463950 642458 463956 642878
rect 464514 642458 464520 642878
rect 463950 642452 464520 642458
rect 464768 642878 465338 642884
rect 464768 642458 464774 642878
rect 465332 642458 465338 642878
rect 462314 641658 462320 642216
rect 462878 641658 462884 642216
rect 464768 642216 465338 642458
rect 465586 642878 466156 643120
rect 465586 642458 465592 642878
rect 466150 642458 466156 642878
rect 465586 642452 466156 642458
rect 466404 642878 466974 643920
rect 468858 644478 469428 644484
rect 468858 643920 468864 644478
rect 469422 643920 469428 644478
rect 466404 642458 466410 642878
rect 466968 642458 466974 642878
rect 466404 642452 466974 642458
rect 467222 642878 467792 642884
rect 467222 642458 467228 642878
rect 467786 642458 467792 642878
rect 468040 642878 468610 642884
rect 468040 642846 468046 642878
rect 468604 642846 468610 642878
rect 468858 642878 469428 643920
rect 471312 644478 471882 644484
rect 471312 643920 471318 644478
rect 471876 643920 471882 644478
rect 464768 641658 464774 642216
rect 465332 641658 465338 642216
rect 467222 642216 467792 642458
rect 467222 641658 467228 642216
rect 467786 641658 467792 642216
rect 467962 642328 467968 642846
rect 468660 642328 468666 642846
rect 468858 642458 468864 642878
rect 469422 642458 469428 642878
rect 468858 642452 469428 642458
rect 469676 643678 470246 643684
rect 469676 643120 469682 643678
rect 470240 643120 470246 643678
rect 469676 642878 470246 643120
rect 469676 642458 469682 642878
rect 470240 642458 470246 642878
rect 469676 642452 470246 642458
rect 470494 642878 471064 642884
rect 470494 642458 470500 642878
rect 471058 642458 471064 642878
rect 462314 641652 462878 641658
rect 464768 641652 465332 641658
rect 467222 641652 467786 641658
rect 467962 641580 468666 642328
rect 470494 642216 471064 642458
rect 471312 642878 471882 643920
rect 473754 642884 474324 646188
rect 482144 646718 482174 646818
rect 482274 646718 482398 646818
rect 482498 646718 482622 646818
rect 482722 646718 482846 646818
rect 482946 646718 483070 646818
rect 483170 646718 483204 646818
rect 482144 646594 483204 646718
rect 482144 646494 482174 646594
rect 482274 646494 482398 646594
rect 482498 646494 482622 646594
rect 482722 646494 482846 646594
rect 482946 646494 483070 646594
rect 483170 646494 483204 646594
rect 482144 646370 483204 646494
rect 482144 646270 482174 646370
rect 482274 646270 482398 646370
rect 482498 646270 482622 646370
rect 482722 646270 482846 646370
rect 482946 646270 483070 646370
rect 483170 646270 483204 646370
rect 482144 646146 483204 646270
rect 482144 646046 482174 646146
rect 482274 646046 482398 646146
rect 482498 646046 482622 646146
rect 482722 646046 482846 646146
rect 482946 646046 483070 646146
rect 483170 646046 483204 646146
rect 482144 645922 483204 646046
rect 482144 645822 482174 645922
rect 482274 645822 482398 645922
rect 482498 645822 482622 645922
rect 482722 645822 482846 645922
rect 482946 645822 483070 645922
rect 483170 645822 483204 645922
rect 482144 645698 483204 645822
rect 482144 645598 482174 645698
rect 482274 645598 482398 645698
rect 482498 645598 482622 645698
rect 482722 645598 482846 645698
rect 482946 645598 483070 645698
rect 483170 645598 483204 645698
rect 482144 645474 483204 645598
rect 482144 645374 482174 645474
rect 482274 645374 482398 645474
rect 482498 645374 482622 645474
rect 482722 645374 482846 645474
rect 482946 645374 483070 645474
rect 483170 645374 483204 645474
rect 482144 645250 483204 645374
rect 482144 645150 482174 645250
rect 482274 645150 482398 645250
rect 482498 645150 482622 645250
rect 482722 645150 482846 645250
rect 482946 645150 483070 645250
rect 483170 645150 483204 645250
rect 482144 645026 483204 645150
rect 482144 644926 482174 645026
rect 482274 644926 482398 645026
rect 482498 644926 482622 645026
rect 482722 644926 482846 645026
rect 482946 644926 483070 645026
rect 483170 644926 483204 645026
rect 482144 644802 483204 644926
rect 482144 644702 482174 644802
rect 482274 644702 482398 644802
rect 482498 644702 482622 644802
rect 482722 644702 482846 644802
rect 482946 644702 483070 644802
rect 483170 644702 483204 644802
rect 482144 644578 483204 644702
rect 482144 644478 482174 644578
rect 482274 644478 482398 644578
rect 482498 644478 482622 644578
rect 482722 644478 482846 644578
rect 482946 644478 483070 644578
rect 483170 644478 483204 644578
rect 482144 644354 483204 644478
rect 482144 644254 482174 644354
rect 482274 644254 482398 644354
rect 482498 644254 482622 644354
rect 482722 644254 482846 644354
rect 482946 644254 483070 644354
rect 483170 644254 483204 644354
rect 482144 644130 483204 644254
rect 482144 644030 482174 644130
rect 482274 644030 482398 644130
rect 482498 644030 482622 644130
rect 482722 644030 482846 644130
rect 482946 644030 483070 644130
rect 483170 644030 483204 644130
rect 482144 643906 483204 644030
rect 482144 643806 482174 643906
rect 482274 643806 482398 643906
rect 482498 643806 482622 643906
rect 482722 643806 482846 643906
rect 482946 643806 483070 643906
rect 483170 643806 483204 643906
rect 482144 643682 483204 643806
rect 482144 643582 482174 643682
rect 482274 643582 482398 643682
rect 482498 643582 482622 643682
rect 482722 643582 482846 643682
rect 482946 643582 483070 643682
rect 483170 643582 483204 643682
rect 482144 643542 483204 643582
rect 471312 642458 471318 642878
rect 471876 642458 471882 642878
rect 471312 642452 471882 642458
rect 472052 642878 472756 642884
rect 470494 641658 470500 642216
rect 471058 641658 471064 642216
rect 472052 642186 472058 642878
rect 472750 642186 472756 642878
rect 472870 642878 473574 642884
rect 472870 642186 472876 642878
rect 473568 642186 473574 642878
rect 473688 642878 474392 642884
rect 473688 642186 473694 642878
rect 474386 642186 474392 642878
rect 472052 642180 472756 642186
rect 473688 642180 474392 642186
rect 470494 641652 471064 641658
rect 459427 641050 459661 641067
rect 459427 640850 459444 641050
rect 459644 640850 459661 641050
rect 459427 640833 459661 640850
rect 459861 641050 460095 641067
rect 459861 640850 459878 641050
rect 460078 640850 460095 641050
rect 459861 640833 460095 640850
rect 460295 641050 460529 641067
rect 460295 640850 460312 641050
rect 460512 640850 460529 641050
rect 460295 640833 460529 640850
rect 460729 641050 460963 641067
rect 460729 640850 460746 641050
rect 460946 640850 460963 641050
rect 460729 640833 460963 640850
rect 461163 641050 461397 641067
rect 461163 640850 461180 641050
rect 461380 640850 461397 641050
rect 461163 640833 461397 640850
rect 461597 641050 461831 641067
rect 461597 640850 461614 641050
rect 461814 640850 461831 641050
rect 461597 640833 461831 640850
rect 462031 641050 462265 641067
rect 462031 640850 462048 641050
rect 462248 640850 462265 641050
rect 462031 640833 462265 640850
rect 462465 641050 462699 641067
rect 462465 640850 462482 641050
rect 462682 640850 462699 641050
rect 462465 640833 462699 640850
rect 462899 641050 463133 641067
rect 462899 640850 462916 641050
rect 463116 640850 463133 641050
rect 462899 640833 463133 640850
rect 463333 641050 463567 641067
rect 463333 640850 463350 641050
rect 463550 640850 463567 641050
rect 463333 640833 463567 640850
rect 463767 641050 464001 641067
rect 463767 640850 463784 641050
rect 463984 640850 464001 641050
rect 463767 640833 464001 640850
rect 464167 641050 464401 641067
rect 464167 640850 464184 641050
rect 464384 640850 464401 641050
rect 464167 640833 464401 640850
rect 464567 641050 464801 641067
rect 464567 640850 464584 641050
rect 464784 640850 464801 641050
rect 464567 640833 464801 640850
rect 464967 641050 465201 641067
rect 464967 640850 464984 641050
rect 465184 640850 465201 641050
rect 464967 640833 465201 640850
rect 465367 641050 465601 641067
rect 465367 640850 465384 641050
rect 465584 640850 465601 641050
rect 465367 640833 465601 640850
rect 465767 641050 466001 641067
rect 465767 640850 465784 641050
rect 465984 640850 466001 641050
rect 465767 640833 466001 640850
rect 466167 641050 466401 641067
rect 466167 640850 466184 641050
rect 466384 640850 466401 641050
rect 466167 640833 466401 640850
rect 466567 641050 466801 641067
rect 466567 640850 466584 641050
rect 466784 640850 466801 641050
rect 466567 640833 466801 640850
rect 466967 641050 467201 641067
rect 466967 640850 466984 641050
rect 467184 640850 467201 641050
rect 466967 640833 467201 640850
rect 467367 641050 467601 641067
rect 467367 640850 467384 641050
rect 467584 640850 467601 641050
rect 467367 640833 467601 640850
rect 459427 640616 459661 640633
rect 459427 640416 459444 640616
rect 459644 640416 459661 640616
rect 459427 640399 459661 640416
rect 459861 640616 460095 640633
rect 459861 640416 459878 640616
rect 460078 640416 460095 640616
rect 459861 640399 460095 640416
rect 460295 640616 460529 640633
rect 460295 640416 460312 640616
rect 460512 640416 460529 640616
rect 460295 640399 460529 640416
rect 460729 640616 460963 640633
rect 460729 640416 460746 640616
rect 460946 640416 460963 640616
rect 460729 640399 460963 640416
rect 461163 640616 461397 640633
rect 461163 640416 461180 640616
rect 461380 640416 461397 640616
rect 461163 640399 461397 640416
rect 461597 640616 461831 640633
rect 461597 640416 461614 640616
rect 461814 640416 461831 640616
rect 461597 640399 461831 640416
rect 462031 640616 462265 640633
rect 462031 640416 462048 640616
rect 462248 640416 462265 640616
rect 462031 640399 462265 640416
rect 462465 640616 462699 640633
rect 462465 640416 462482 640616
rect 462682 640416 462699 640616
rect 462465 640399 462699 640416
rect 462899 640616 463133 640633
rect 462899 640416 462916 640616
rect 463116 640416 463133 640616
rect 462899 640399 463133 640416
rect 463333 640616 463567 640633
rect 463333 640416 463350 640616
rect 463550 640416 463567 640616
rect 463333 640399 463567 640416
rect 463767 640616 464001 640633
rect 463767 640416 463784 640616
rect 463984 640416 464001 640616
rect 463767 640399 464001 640416
rect 467962 640334 468664 641580
rect 468967 641050 469201 641067
rect 468967 640850 468984 641050
rect 469184 640850 469201 641050
rect 468967 640833 469201 640850
rect 469367 641050 469601 641067
rect 469367 640850 469384 641050
rect 469584 640850 469601 641050
rect 469367 640833 469601 640850
rect 469767 641050 470001 641067
rect 469767 640850 469784 641050
rect 469984 640850 470001 641050
rect 469767 640833 470001 640850
rect 470167 641050 470401 641067
rect 470167 640850 470184 641050
rect 470384 640850 470401 641050
rect 470167 640833 470401 640850
rect 470567 641050 470801 641067
rect 470567 640850 470584 641050
rect 470784 640850 470801 641050
rect 470567 640833 470801 640850
rect 470967 641050 471201 641067
rect 470967 640850 470984 641050
rect 471184 640850 471201 641050
rect 470967 640833 471201 640850
rect 471367 641050 471601 641067
rect 471367 640850 471384 641050
rect 471584 640850 471601 641050
rect 471367 640833 471601 640850
rect 471767 641050 472001 641067
rect 471767 640850 471784 641050
rect 471984 640850 472001 641050
rect 471767 640833 472001 640850
rect 472167 641050 472401 641067
rect 472167 640850 472184 641050
rect 472384 640850 472401 641050
rect 472167 640833 472401 640850
rect 467962 640328 472474 640334
rect 459427 640182 459661 640199
rect 459427 639982 459444 640182
rect 459644 639982 459661 640182
rect 459427 639965 459661 639982
rect 459861 640182 460095 640199
rect 459861 639982 459878 640182
rect 460078 639982 460095 640182
rect 459861 639965 460095 639982
rect 460295 640182 460529 640199
rect 460295 639982 460312 640182
rect 460512 639982 460529 640182
rect 460295 639965 460529 639982
rect 460729 640182 460963 640199
rect 460729 639982 460746 640182
rect 460946 639982 460963 640182
rect 460729 639965 460963 639982
rect 461163 640182 461397 640199
rect 461163 639982 461180 640182
rect 461380 639982 461397 640182
rect 461163 639965 461397 639982
rect 461597 640182 461831 640199
rect 461597 639982 461614 640182
rect 461814 639982 461831 640182
rect 461597 639965 461831 639982
rect 462031 640182 462265 640199
rect 462031 639982 462048 640182
rect 462248 639982 462265 640182
rect 462031 639965 462265 639982
rect 462465 640182 462699 640199
rect 462465 639982 462482 640182
rect 462682 639982 462699 640182
rect 462465 639965 462699 639982
rect 462899 640182 463133 640199
rect 462899 639982 462916 640182
rect 463116 639982 463133 640182
rect 462899 639965 463133 639982
rect 463333 640182 463567 640199
rect 463333 639982 463350 640182
rect 463550 639982 463567 640182
rect 463333 639965 463567 639982
rect 463767 640182 464001 640199
rect 463767 639982 463784 640182
rect 463984 639982 464001 640182
rect 463767 639965 464001 639982
rect 467962 639810 471534 640328
rect 472468 639810 472474 640328
rect 467962 639804 472474 639810
rect 452342 639548 473588 639556
rect 452342 639474 453864 639548
rect 455852 639474 467564 639548
rect 469552 639474 472876 639548
rect 452342 638798 452996 639474
rect 473568 639098 473588 639548
rect 452340 638792 452996 638798
rect 452340 638378 452346 638792
rect 452466 638490 452996 638792
rect 473318 638490 473588 639098
rect 452466 638396 453864 638490
rect 455852 638396 467564 638490
rect 469552 638396 473588 638490
rect 452466 638378 473588 638396
rect 452340 638374 473588 638378
rect 452340 638372 452472 638374
rect 443004 638212 443594 638272
rect 443004 638152 443024 638212
rect 443084 638152 443144 638212
rect 443204 638152 443264 638212
rect 443324 638152 443384 638212
rect 443444 638152 443504 638212
rect 443564 638152 443594 638212
rect 443004 638092 443594 638152
rect 443004 638032 443024 638092
rect 443084 638032 443144 638092
rect 443204 638032 443264 638092
rect 443324 638032 443384 638092
rect 443444 638032 443504 638092
rect 443564 638032 443594 638092
rect 437864 636778 438922 636788
rect 437864 636678 437894 636778
rect 437994 636678 438118 636778
rect 438218 636678 438342 636778
rect 438442 636678 438566 636778
rect 438666 636678 438790 636778
rect 438890 636678 438922 636778
rect 437864 636554 438922 636678
rect 437864 636454 437894 636554
rect 437994 636454 438118 636554
rect 438218 636454 438342 636554
rect 438442 636454 438566 636554
rect 438666 636454 438790 636554
rect 438890 636454 438922 636554
rect 437864 636330 438922 636454
rect 437864 636230 437894 636330
rect 437994 636230 438118 636330
rect 438218 636230 438342 636330
rect 438442 636230 438566 636330
rect 438666 636230 438790 636330
rect 438890 636230 438922 636330
rect 437864 636106 438922 636230
rect 443004 636366 443594 638032
rect 451884 638086 474392 638090
rect 451884 637794 451890 638086
rect 452010 638084 474392 638086
rect 452010 637796 456564 638084
rect 458552 637796 464864 638084
rect 466852 637796 473696 638084
rect 474386 637796 474392 638084
rect 452010 637794 474392 637796
rect 451884 637490 474392 637794
rect 443004 636296 443016 636366
rect 443076 636296 443088 636366
rect 443148 636296 443160 636366
rect 443220 636296 443232 636366
rect 443292 636296 443304 636366
rect 443364 636296 443376 636366
rect 443436 636296 443448 636366
rect 443508 636296 443520 636366
rect 443580 636296 443594 636366
rect 443004 636272 443594 636296
rect 443004 636202 443016 636272
rect 443076 636202 443088 636272
rect 443148 636202 443160 636272
rect 443220 636202 443232 636272
rect 443292 636202 443304 636272
rect 443364 636202 443376 636272
rect 443436 636202 443448 636272
rect 443508 636202 443520 636272
rect 443580 636202 443594 636272
rect 443004 636192 443594 636202
rect 482144 636778 483202 636788
rect 482144 636678 482174 636778
rect 482274 636678 482398 636778
rect 482498 636678 482622 636778
rect 482722 636678 482846 636778
rect 482946 636678 483070 636778
rect 483170 636678 483202 636778
rect 482144 636554 483202 636678
rect 482144 636454 482174 636554
rect 482274 636454 482398 636554
rect 482498 636454 482622 636554
rect 482722 636454 482846 636554
rect 482946 636454 483070 636554
rect 483170 636454 483202 636554
rect 482144 636330 483202 636454
rect 482144 636230 482174 636330
rect 482274 636230 482398 636330
rect 482498 636230 482622 636330
rect 482722 636230 482846 636330
rect 482946 636230 483070 636330
rect 483170 636230 483202 636330
rect 437864 636006 437894 636106
rect 437994 636006 438118 636106
rect 438218 636006 438342 636106
rect 438442 636006 438566 636106
rect 438666 636006 438790 636106
rect 438890 636006 438922 636106
rect 437864 635882 438922 636006
rect 437864 635782 437894 635882
rect 437994 635782 438118 635882
rect 438218 635782 438342 635882
rect 438442 635782 438566 635882
rect 438666 635782 438790 635882
rect 438890 635782 438922 635882
rect 437864 635658 438922 635782
rect 482144 636106 483202 636230
rect 482144 636006 482174 636106
rect 482274 636006 482398 636106
rect 482498 636006 482622 636106
rect 482722 636006 482846 636106
rect 482946 636006 483070 636106
rect 483170 636006 483202 636106
rect 482144 635882 483202 636006
rect 482144 635782 482174 635882
rect 482274 635782 482398 635882
rect 482498 635782 482622 635882
rect 482722 635782 482846 635882
rect 482946 635782 483070 635882
rect 483170 635782 483202 635882
rect 437864 635558 437894 635658
rect 437994 635558 438118 635658
rect 438218 635558 438342 635658
rect 438442 635558 438566 635658
rect 438666 635558 438790 635658
rect 438890 635558 438922 635658
rect 437864 635434 438922 635558
rect 437864 635334 437894 635434
rect 437994 635334 438118 635434
rect 438218 635334 438342 635434
rect 438442 635334 438566 635434
rect 438666 635334 438790 635434
rect 438890 635334 438922 635434
rect 437864 635210 438922 635334
rect 437864 635110 437894 635210
rect 437994 635110 438118 635210
rect 438218 635110 438342 635210
rect 438442 635110 438566 635210
rect 438666 635110 438790 635210
rect 438890 635110 438922 635210
rect 437864 634986 438922 635110
rect 472870 635760 478264 635766
rect 472870 635068 472876 635760
rect 473568 635702 478264 635760
rect 473568 635650 477640 635702
rect 477692 635650 477744 635702
rect 477796 635650 477848 635702
rect 477900 635650 477952 635702
rect 478004 635650 478056 635702
rect 478108 635650 478160 635702
rect 478212 635650 478264 635702
rect 473568 635598 478264 635650
rect 473568 635546 477640 635598
rect 477692 635546 477744 635598
rect 477796 635546 477848 635598
rect 477900 635546 477952 635598
rect 478004 635546 478056 635598
rect 478108 635546 478160 635598
rect 478212 635546 478264 635598
rect 473568 635494 478264 635546
rect 473568 635442 477640 635494
rect 477692 635442 477744 635494
rect 477796 635442 477848 635494
rect 477900 635442 477952 635494
rect 478004 635442 478056 635494
rect 478108 635442 478160 635494
rect 478212 635442 478264 635494
rect 473568 635390 478264 635442
rect 473568 635338 477640 635390
rect 477692 635338 477744 635390
rect 477796 635338 477848 635390
rect 477900 635338 477952 635390
rect 478004 635338 478056 635390
rect 478108 635338 478160 635390
rect 478212 635338 478264 635390
rect 473568 635286 478264 635338
rect 473568 635234 477640 635286
rect 477692 635234 477744 635286
rect 477796 635234 477848 635286
rect 477900 635234 477952 635286
rect 478004 635234 478056 635286
rect 478108 635234 478160 635286
rect 478212 635234 478264 635286
rect 473568 635182 478264 635234
rect 473568 635130 477640 635182
rect 477692 635130 477744 635182
rect 477796 635130 477848 635182
rect 477900 635130 477952 635182
rect 478004 635130 478056 635182
rect 478108 635130 478160 635182
rect 478212 635130 478264 635182
rect 473568 635068 478264 635130
rect 472870 635062 478264 635068
rect 482144 635658 483202 635782
rect 482144 635558 482174 635658
rect 482274 635558 482398 635658
rect 482498 635558 482622 635658
rect 482722 635558 482846 635658
rect 482946 635558 483070 635658
rect 483170 635558 483202 635658
rect 482144 635434 483202 635558
rect 482144 635334 482174 635434
rect 482274 635334 482398 635434
rect 482498 635334 482622 635434
rect 482722 635334 482846 635434
rect 482946 635334 483070 635434
rect 483170 635334 483202 635434
rect 482144 635210 483202 635334
rect 482144 635110 482174 635210
rect 482274 635110 482398 635210
rect 482498 635110 482622 635210
rect 482722 635110 482846 635210
rect 482946 635110 483070 635210
rect 483170 635110 483202 635210
rect 437864 634886 437894 634986
rect 437994 634886 438118 634986
rect 438218 634886 438342 634986
rect 438442 634886 438566 634986
rect 438666 634886 438790 634986
rect 438890 634886 438922 634986
rect 437864 634762 438922 634886
rect 437864 634662 437894 634762
rect 437994 634662 438118 634762
rect 438218 634662 438342 634762
rect 438442 634662 438566 634762
rect 438666 634662 438790 634762
rect 438890 634662 438922 634762
rect 482144 634986 483202 635110
rect 482144 634886 482174 634986
rect 482274 634886 482398 634986
rect 482498 634886 482622 634986
rect 482722 634886 482846 634986
rect 482946 634886 483070 634986
rect 483170 634886 483202 634986
rect 482144 634762 483202 634886
rect 437864 634538 438922 634662
rect 446664 634674 452346 634694
rect 446664 634620 446684 634674
rect 446828 634620 447828 634674
rect 447972 634620 448972 634674
rect 449116 634620 452346 634674
rect 446664 634614 452346 634620
rect 452466 634614 452472 634694
rect 482144 634662 482174 634762
rect 482274 634662 482398 634762
rect 482498 634662 482622 634762
rect 482722 634662 482846 634762
rect 482946 634662 483070 634762
rect 483170 634662 483202 634762
rect 437864 634438 437894 634538
rect 437994 634438 438118 634538
rect 438218 634438 438342 634538
rect 438442 634438 438566 634538
rect 438666 634438 438790 634538
rect 438890 634438 438922 634538
rect 446092 634534 451890 634554
rect 446092 634480 446112 634534
rect 446256 634480 447256 634534
rect 447400 634480 448400 634534
rect 448544 634480 451890 634534
rect 446092 634474 451890 634480
rect 452000 634474 452006 634554
rect 482144 634538 483202 634662
rect 437864 634314 438922 634438
rect 437864 634214 437894 634314
rect 437994 634214 438118 634314
rect 438218 634214 438342 634314
rect 438442 634214 438566 634314
rect 438666 634214 438790 634314
rect 438890 634214 438922 634314
rect 437864 634090 438922 634214
rect 437864 633990 437894 634090
rect 437994 633990 438118 634090
rect 438218 633990 438342 634090
rect 438442 633990 438566 634090
rect 438666 633990 438790 634090
rect 438890 633990 438922 634090
rect 437864 633866 438922 633990
rect 437864 633766 437894 633866
rect 437994 633766 438118 633866
rect 438218 633766 438342 633866
rect 438442 633766 438566 633866
rect 438666 633766 438790 633866
rect 438890 633766 438922 633866
rect 437864 633642 438922 633766
rect 437864 633542 437894 633642
rect 437994 633542 438118 633642
rect 438218 633542 438342 633642
rect 438442 633542 438566 633642
rect 438666 633542 438790 633642
rect 438890 633542 438922 633642
rect 437864 633418 438922 633542
rect 437864 633318 437894 633418
rect 437994 633318 438118 633418
rect 438218 633318 438342 633418
rect 438442 633318 438566 633418
rect 438666 633318 438790 633418
rect 438890 633318 438922 633418
rect 437864 633194 438922 633318
rect 437864 633094 437894 633194
rect 437994 633094 438118 633194
rect 438218 633094 438342 633194
rect 438442 633094 438566 633194
rect 438666 633094 438790 633194
rect 438890 633094 438922 633194
rect 437864 632970 438922 633094
rect 437864 632870 437894 632970
rect 437994 632870 438118 632970
rect 438218 632870 438342 632970
rect 438442 632870 438566 632970
rect 438666 632870 438790 632970
rect 438890 632870 438922 632970
rect 437864 632746 438922 632870
rect 437864 632646 437894 632746
rect 437994 632646 438118 632746
rect 438218 632646 438342 632746
rect 438442 632646 438566 632746
rect 438666 632646 438790 632746
rect 438890 632646 438922 632746
rect 482144 634438 482174 634538
rect 482274 634438 482398 634538
rect 482498 634438 482622 634538
rect 482722 634438 482846 634538
rect 482946 634438 483070 634538
rect 483170 634438 483202 634538
rect 482144 634314 483202 634438
rect 482144 634214 482174 634314
rect 482274 634214 482398 634314
rect 482498 634214 482622 634314
rect 482722 634214 482846 634314
rect 482946 634214 483070 634314
rect 483170 634214 483202 634314
rect 482144 634090 483202 634214
rect 482144 633990 482174 634090
rect 482274 633990 482398 634090
rect 482498 633990 482622 634090
rect 482722 633990 482846 634090
rect 482946 633990 483070 634090
rect 483170 633990 483202 634090
rect 482144 633866 483202 633990
rect 482144 633766 482174 633866
rect 482274 633766 482398 633866
rect 482498 633766 482622 633866
rect 482722 633766 482846 633866
rect 482946 633766 483070 633866
rect 483170 633766 483202 633866
rect 482144 633642 483202 633766
rect 482144 633542 482174 633642
rect 482274 633542 482398 633642
rect 482498 633542 482622 633642
rect 482722 633542 482846 633642
rect 482946 633542 483070 633642
rect 483170 633542 483202 633642
rect 482144 633418 483202 633542
rect 482144 633318 482174 633418
rect 482274 633318 482398 633418
rect 482498 633318 482622 633418
rect 482722 633318 482846 633418
rect 482946 633318 483070 633418
rect 483170 633318 483202 633418
rect 482144 633194 483202 633318
rect 482144 633094 482174 633194
rect 482274 633094 482398 633194
rect 482498 633094 482622 633194
rect 482722 633094 482846 633194
rect 482946 633094 483070 633194
rect 483170 633094 483202 633194
rect 482144 632970 483202 633094
rect 482144 632870 482174 632970
rect 482274 632870 482398 632970
rect 482498 632870 482622 632970
rect 482722 632870 482846 632970
rect 482946 632870 483070 632970
rect 483170 632870 483202 632970
rect 482144 632746 483202 632870
rect 437864 632522 438922 632646
rect 440878 632690 443524 632696
rect 440878 632684 442718 632690
rect 440878 632632 440884 632684
rect 440936 632638 442718 632684
rect 442770 632638 443324 632690
rect 440936 632632 443324 632638
rect 443518 632632 443524 632690
rect 440878 632626 443524 632632
rect 482144 632646 482174 632746
rect 482274 632646 482398 632746
rect 482498 632646 482622 632746
rect 482722 632646 482846 632746
rect 482946 632646 483070 632746
rect 483170 632646 483202 632746
rect 437864 632422 437894 632522
rect 437994 632422 438118 632522
rect 438218 632422 438342 632522
rect 438442 632422 438566 632522
rect 438666 632422 438790 632522
rect 438890 632422 438922 632522
rect 482144 632522 483202 632646
rect 437864 632298 438922 632422
rect 440931 632478 449302 632486
rect 440931 632426 441802 632478
rect 441854 632468 449302 632478
rect 441854 632426 446380 632468
rect 440931 632364 446380 632426
rect 446432 632364 446952 632468
rect 447004 632364 447524 632468
rect 447576 632364 448096 632468
rect 448148 632364 448668 632468
rect 448720 632364 449240 632468
rect 449292 632364 449302 632468
rect 440931 632352 449302 632364
rect 482144 632422 482174 632522
rect 482274 632422 482398 632522
rect 482498 632422 482622 632522
rect 482722 632422 482846 632522
rect 482946 632422 483070 632522
rect 483170 632422 483202 632522
rect 437864 632198 437894 632298
rect 437994 632198 438118 632298
rect 438218 632198 438342 632298
rect 438442 632198 438566 632298
rect 438666 632198 438790 632298
rect 438890 632198 438922 632298
rect 437864 632074 438922 632198
rect 437864 631974 437894 632074
rect 437994 631974 438118 632074
rect 438218 631974 438342 632074
rect 438442 631974 438566 632074
rect 438666 631974 438790 632074
rect 438890 631974 438922 632074
rect 443628 632318 453232 632324
rect 443628 632317 444480 632318
rect 443628 632065 443648 632317
rect 444248 632065 444480 632317
rect 443628 632064 444480 632065
rect 444532 632064 445040 632318
rect 445092 632064 445600 632318
rect 445652 632064 446500 632318
rect 446552 632064 447644 632318
rect 447696 632064 448788 632318
rect 448840 632064 449588 632318
rect 449640 632064 450148 632318
rect 450200 632064 450708 632318
rect 450760 632317 452758 632318
rect 450760 632065 452139 632317
rect 452739 632065 452758 632317
rect 450760 632064 452758 632065
rect 453226 632064 453232 632318
rect 443628 632058 453232 632064
rect 482144 632298 483202 632422
rect 482144 632198 482174 632298
rect 482274 632198 482398 632298
rect 482498 632198 482622 632298
rect 482722 632198 482846 632298
rect 482946 632198 483070 632298
rect 483170 632198 483202 632298
rect 482144 632074 483202 632198
rect 437864 631850 438922 631974
rect 446072 632028 449152 632030
rect 446072 631970 446078 632028
rect 446286 632024 447222 632028
rect 446286 631970 446650 632024
rect 446072 631966 446650 631970
rect 446858 631970 447222 632024
rect 447430 631970 447794 632028
rect 448002 631970 448366 632028
rect 448574 631970 448938 632028
rect 449146 631970 449152 632028
rect 446858 631966 449152 631970
rect 446072 631964 449152 631966
rect 482144 631974 482174 632074
rect 482274 631974 482398 632074
rect 482498 631974 482622 632074
rect 482722 631974 482846 632074
rect 482946 631974 483070 632074
rect 483170 631974 483202 632074
rect 446072 631960 447118 631964
rect 437864 631750 437894 631850
rect 437994 631750 438118 631850
rect 438218 631750 438342 631850
rect 438442 631750 438566 631850
rect 438666 631750 438790 631850
rect 438890 631750 438922 631850
rect 437864 631626 438922 631750
rect 437864 631526 437894 631626
rect 437994 631526 438118 631626
rect 438218 631526 438342 631626
rect 438442 631526 438566 631626
rect 438666 631526 438790 631626
rect 438890 631526 438922 631626
rect 437864 631402 438922 631526
rect 437864 631302 437894 631402
rect 437994 631302 438118 631402
rect 438218 631302 438342 631402
rect 438442 631302 438566 631402
rect 438666 631302 438790 631402
rect 438890 631302 438922 631402
rect 437864 631178 438922 631302
rect 437864 631078 437894 631178
rect 437994 631078 438118 631178
rect 438218 631078 438342 631178
rect 438442 631078 438566 631178
rect 438666 631078 438790 631178
rect 438890 631078 438922 631178
rect 437864 630954 438922 631078
rect 437864 630854 437894 630954
rect 437994 630854 438118 630954
rect 438218 630854 438342 630954
rect 438442 630854 438566 630954
rect 438666 630854 438790 630954
rect 438890 630854 438922 630954
rect 482144 631850 483202 631974
rect 482144 631750 482174 631850
rect 482274 631750 482398 631850
rect 482498 631750 482622 631850
rect 482722 631750 482846 631850
rect 482946 631750 483070 631850
rect 483170 631750 483202 631850
rect 482144 631626 483202 631750
rect 482144 631526 482174 631626
rect 482274 631526 482398 631626
rect 482498 631526 482622 631626
rect 482722 631526 482846 631626
rect 482946 631526 483070 631626
rect 483170 631526 483202 631626
rect 482144 631402 483202 631526
rect 482144 631302 482174 631402
rect 482274 631302 482398 631402
rect 482498 631302 482622 631402
rect 482722 631302 482846 631402
rect 482946 631302 483070 631402
rect 483170 631302 483202 631402
rect 482144 631178 483202 631302
rect 482144 631078 482174 631178
rect 482274 631078 482398 631178
rect 482498 631078 482622 631178
rect 482722 631078 482846 631178
rect 482946 631078 483070 631178
rect 483170 631078 483202 631178
rect 482144 630954 483202 631078
rect 437864 630730 438922 630854
rect 437864 630630 437894 630730
rect 437994 630630 438118 630730
rect 438218 630630 438342 630730
rect 438442 630630 438566 630730
rect 438666 630630 438790 630730
rect 438890 630630 438922 630730
rect 437864 630506 438922 630630
rect 437864 630406 437894 630506
rect 437994 630406 438118 630506
rect 438218 630406 438342 630506
rect 438442 630406 438566 630506
rect 438666 630406 438790 630506
rect 438890 630406 438922 630506
rect 437864 630282 438922 630406
rect 437864 630182 437894 630282
rect 437994 630182 438118 630282
rect 438218 630182 438342 630282
rect 438442 630182 438566 630282
rect 438666 630182 438790 630282
rect 438890 630182 438922 630282
rect 437864 630162 438922 630182
rect 471526 630850 477016 630856
rect 471526 629914 471532 630850
rect 472468 630550 477016 630850
rect 472468 630498 476352 630550
rect 476404 630498 476456 630550
rect 476508 630498 476560 630550
rect 476612 630498 476664 630550
rect 476716 630498 476768 630550
rect 476820 630498 476872 630550
rect 476924 630498 477016 630550
rect 472468 630446 477016 630498
rect 472468 630394 476352 630446
rect 476404 630394 476456 630446
rect 476508 630394 476560 630446
rect 476612 630394 476664 630446
rect 476716 630394 476768 630446
rect 476820 630394 476872 630446
rect 476924 630394 477016 630446
rect 472468 630342 477016 630394
rect 472468 630290 476352 630342
rect 476404 630290 476456 630342
rect 476508 630290 476560 630342
rect 476612 630290 476664 630342
rect 476716 630290 476768 630342
rect 476820 630290 476872 630342
rect 476924 630290 477016 630342
rect 472468 630238 477016 630290
rect 472468 630186 476352 630238
rect 476404 630186 476456 630238
rect 476508 630186 476560 630238
rect 476612 630186 476664 630238
rect 476716 630186 476768 630238
rect 476820 630186 476872 630238
rect 476924 630186 477016 630238
rect 472468 630134 477016 630186
rect 482144 630854 482174 630954
rect 482274 630854 482398 630954
rect 482498 630854 482622 630954
rect 482722 630854 482846 630954
rect 482946 630854 483070 630954
rect 483170 630854 483202 630954
rect 482144 630730 483202 630854
rect 482144 630630 482174 630730
rect 482274 630630 482398 630730
rect 482498 630630 482622 630730
rect 482722 630630 482846 630730
rect 482946 630630 483070 630730
rect 483170 630630 483202 630730
rect 482144 630506 483202 630630
rect 482144 630406 482174 630506
rect 482274 630406 482398 630506
rect 482498 630406 482622 630506
rect 482722 630406 482846 630506
rect 482946 630406 483070 630506
rect 483170 630406 483202 630506
rect 482144 630282 483202 630406
rect 482144 630182 482174 630282
rect 482274 630182 482398 630282
rect 482498 630182 482622 630282
rect 482722 630182 482846 630282
rect 482946 630182 483070 630282
rect 483170 630182 483202 630282
rect 482144 630162 483202 630182
rect 472468 630082 476352 630134
rect 476404 630082 476456 630134
rect 476508 630082 476560 630134
rect 476612 630082 476664 630134
rect 476716 630082 476768 630134
rect 476820 630082 476872 630134
rect 476924 630082 477016 630134
rect 472468 630030 477016 630082
rect 472468 629978 476352 630030
rect 476404 629978 476456 630030
rect 476508 629978 476560 630030
rect 476612 629978 476664 630030
rect 476716 629978 476768 630030
rect 476820 629978 476872 630030
rect 476924 629978 477016 630030
rect 472468 629914 477016 629978
rect 471526 629908 477016 629914
rect 442980 629244 452246 629250
rect 442980 629130 442990 629244
rect 452236 629130 452246 629244
rect 442980 629126 452246 629130
rect 452752 629224 469378 629230
rect 452752 629076 452758 629224
rect 453226 629210 469378 629224
rect 453226 629090 454078 629210
rect 454218 629090 454538 629210
rect 454678 629090 454998 629210
rect 455138 629090 455458 629210
rect 455598 629090 455918 629210
rect 456058 629090 456378 629210
rect 456518 629090 456838 629210
rect 456978 629090 457298 629210
rect 457438 629090 457758 629210
rect 457898 629090 458218 629210
rect 458358 629090 459578 629210
rect 459718 629090 460038 629210
rect 460178 629090 460498 629210
rect 460638 629090 460958 629210
rect 461098 629090 461418 629210
rect 461558 629090 461878 629210
rect 462018 629090 462338 629210
rect 462478 629090 462798 629210
rect 462938 629090 463258 629210
rect 463398 629090 463718 629210
rect 463858 629090 465078 629210
rect 465218 629090 465538 629210
rect 465678 629090 465998 629210
rect 466138 629090 466458 629210
rect 466598 629090 466918 629210
rect 467058 629090 467378 629210
rect 467518 629090 467838 629210
rect 467978 629090 468298 629210
rect 468438 629090 468758 629210
rect 468898 629090 469218 629210
rect 469358 629090 469378 629210
rect 453226 629076 469378 629090
rect 452752 629070 469378 629076
rect 443318 629050 443524 629052
rect 443318 629046 450558 629050
rect 443318 628932 443324 629046
rect 443518 629040 450558 629046
rect 443518 628936 444204 629040
rect 444256 628936 444776 629040
rect 444828 628936 445348 629040
rect 445400 628936 449352 629040
rect 449404 628936 449924 629040
rect 449976 628936 450496 629040
rect 450548 628936 450558 629040
rect 454318 629022 454438 629030
rect 455238 629022 455358 629030
rect 456158 629022 456278 629030
rect 457078 629022 457198 629030
rect 457998 629022 458118 629030
rect 459818 629022 459938 629030
rect 460738 629022 460858 629030
rect 461658 629022 461778 629030
rect 462578 629022 462698 629030
rect 463498 629022 463618 629030
rect 465318 629022 465438 629030
rect 466238 629022 466358 629030
rect 467158 629022 467278 629030
rect 468078 629022 468198 629030
rect 468998 629022 469118 629030
rect 443518 628932 450558 628936
rect 443318 628926 450558 628932
rect 452744 629012 470702 629022
rect 452744 628694 452754 629012
rect 470692 628988 470702 629012
rect 470692 628694 470714 628988
rect 452744 628688 470714 628694
rect 452744 628686 470702 628688
rect 438880 627656 445540 627686
rect 438880 627556 438920 627656
rect 439020 627556 439144 627656
rect 439244 627556 439368 627656
rect 439468 627556 439592 627656
rect 439692 627556 439816 627656
rect 439916 627556 440040 627656
rect 440140 627556 440264 627656
rect 440364 627556 440488 627656
rect 440588 627556 440712 627656
rect 440812 627556 440936 627656
rect 441036 627556 441160 627656
rect 441260 627556 441384 627656
rect 441484 627556 441608 627656
rect 441708 627556 441832 627656
rect 441932 627556 442056 627656
rect 442156 627556 442280 627656
rect 442380 627556 442504 627656
rect 442604 627556 442728 627656
rect 442828 627556 442952 627656
rect 443052 627556 443176 627656
rect 443276 627556 443400 627656
rect 443500 627556 443624 627656
rect 443724 627556 443848 627656
rect 443948 627556 444072 627656
rect 444172 627556 444296 627656
rect 444396 627556 444520 627656
rect 444620 627556 444744 627656
rect 444844 627556 444968 627656
rect 445068 627556 445192 627656
rect 445292 627556 445416 627656
rect 445516 627556 445540 627656
rect 438880 627432 445540 627556
rect 438880 627332 438920 627432
rect 439020 627332 439144 627432
rect 439244 627332 439368 627432
rect 439468 627332 439592 627432
rect 439692 627332 439816 627432
rect 439916 627332 440040 627432
rect 440140 627332 440264 627432
rect 440364 627332 440488 627432
rect 440588 627332 440712 627432
rect 440812 627332 440936 627432
rect 441036 627332 441160 627432
rect 441260 627332 441384 627432
rect 441484 627332 441608 627432
rect 441708 627332 441832 627432
rect 441932 627332 442056 627432
rect 442156 627332 442280 627432
rect 442380 627332 442504 627432
rect 442604 627332 442728 627432
rect 442828 627332 442952 627432
rect 443052 627332 443176 627432
rect 443276 627332 443400 627432
rect 443500 627332 443624 627432
rect 443724 627332 443848 627432
rect 443948 627332 444072 627432
rect 444172 627332 444296 627432
rect 444396 627332 444520 627432
rect 444620 627332 444744 627432
rect 444844 627332 444968 627432
rect 445068 627332 445192 627432
rect 445292 627332 445416 627432
rect 445516 627332 445540 627432
rect 438880 627208 445540 627332
rect 438880 627108 438920 627208
rect 439020 627108 439144 627208
rect 439244 627108 439368 627208
rect 439468 627108 439592 627208
rect 439692 627108 439816 627208
rect 439916 627108 440040 627208
rect 440140 627108 440264 627208
rect 440364 627108 440488 627208
rect 440588 627108 440712 627208
rect 440812 627108 440936 627208
rect 441036 627108 441160 627208
rect 441260 627108 441384 627208
rect 441484 627108 441608 627208
rect 441708 627108 441832 627208
rect 441932 627108 442056 627208
rect 442156 627108 442280 627208
rect 442380 627108 442504 627208
rect 442604 627108 442728 627208
rect 442828 627108 442952 627208
rect 443052 627108 443176 627208
rect 443276 627108 443400 627208
rect 443500 627108 443624 627208
rect 443724 627108 443848 627208
rect 443948 627108 444072 627208
rect 444172 627108 444296 627208
rect 444396 627108 444520 627208
rect 444620 627108 444744 627208
rect 444844 627108 444968 627208
rect 445068 627108 445192 627208
rect 445292 627108 445416 627208
rect 445516 627108 445540 627208
rect 438880 626984 445540 627108
rect 438880 626884 438920 626984
rect 439020 626884 439144 626984
rect 439244 626884 439368 626984
rect 439468 626884 439592 626984
rect 439692 626884 439816 626984
rect 439916 626884 440040 626984
rect 440140 626884 440264 626984
rect 440364 626884 440488 626984
rect 440588 626884 440712 626984
rect 440812 626884 440936 626984
rect 441036 626884 441160 626984
rect 441260 626884 441384 626984
rect 441484 626884 441608 626984
rect 441708 626884 441832 626984
rect 441932 626884 442056 626984
rect 442156 626884 442280 626984
rect 442380 626884 442504 626984
rect 442604 626884 442728 626984
rect 442828 626884 442952 626984
rect 443052 626884 443176 626984
rect 443276 626884 443400 626984
rect 443500 626884 443624 626984
rect 443724 626884 443848 626984
rect 443948 626884 444072 626984
rect 444172 626884 444296 626984
rect 444396 626884 444520 626984
rect 444620 626884 444744 626984
rect 444844 626884 444968 626984
rect 445068 626884 445192 626984
rect 445292 626884 445416 626984
rect 445516 626884 445540 626984
rect 438880 626760 445540 626884
rect 438880 626660 438920 626760
rect 439020 626660 439144 626760
rect 439244 626660 439368 626760
rect 439468 626660 439592 626760
rect 439692 626660 439816 626760
rect 439916 626660 440040 626760
rect 440140 626660 440264 626760
rect 440364 626660 440488 626760
rect 440588 626660 440712 626760
rect 440812 626660 440936 626760
rect 441036 626660 441160 626760
rect 441260 626660 441384 626760
rect 441484 626660 441608 626760
rect 441708 626660 441832 626760
rect 441932 626660 442056 626760
rect 442156 626660 442280 626760
rect 442380 626660 442504 626760
rect 442604 626660 442728 626760
rect 442828 626660 442952 626760
rect 443052 626660 443176 626760
rect 443276 626660 443400 626760
rect 443500 626660 443624 626760
rect 443724 626660 443848 626760
rect 443948 626660 444072 626760
rect 444172 626660 444296 626760
rect 444396 626660 444520 626760
rect 444620 626660 444744 626760
rect 444844 626660 444968 626760
rect 445068 626660 445192 626760
rect 445292 626660 445416 626760
rect 445516 626660 445540 626760
rect 438880 626626 445540 626660
rect 449350 627656 456010 627686
rect 449350 627556 449390 627656
rect 449490 627556 449614 627656
rect 449714 627556 449838 627656
rect 449938 627556 450062 627656
rect 450162 627556 450286 627656
rect 450386 627556 450510 627656
rect 450610 627556 450734 627656
rect 450834 627556 450958 627656
rect 451058 627556 451182 627656
rect 451282 627556 451406 627656
rect 451506 627556 451630 627656
rect 451730 627556 451854 627656
rect 451954 627556 452078 627656
rect 452178 627556 452302 627656
rect 452402 627556 452526 627656
rect 452626 627556 452750 627656
rect 452850 627556 452974 627656
rect 453074 627556 453198 627656
rect 453298 627556 453422 627656
rect 453522 627556 453646 627656
rect 453746 627556 453870 627656
rect 453970 627556 454094 627656
rect 454194 627556 454318 627656
rect 454418 627556 454542 627656
rect 454642 627556 454766 627656
rect 454866 627556 454990 627656
rect 455090 627556 455214 627656
rect 455314 627556 455438 627656
rect 455538 627556 455662 627656
rect 455762 627556 455886 627656
rect 455986 627556 456010 627656
rect 449350 627432 456010 627556
rect 449350 627332 449390 627432
rect 449490 627332 449614 627432
rect 449714 627332 449838 627432
rect 449938 627332 450062 627432
rect 450162 627332 450286 627432
rect 450386 627332 450510 627432
rect 450610 627332 450734 627432
rect 450834 627332 450958 627432
rect 451058 627332 451182 627432
rect 451282 627332 451406 627432
rect 451506 627332 451630 627432
rect 451730 627332 451854 627432
rect 451954 627332 452078 627432
rect 452178 627332 452302 627432
rect 452402 627332 452526 627432
rect 452626 627332 452750 627432
rect 452850 627332 452974 627432
rect 453074 627332 453198 627432
rect 453298 627332 453422 627432
rect 453522 627332 453646 627432
rect 453746 627332 453870 627432
rect 453970 627332 454094 627432
rect 454194 627332 454318 627432
rect 454418 627332 454542 627432
rect 454642 627332 454766 627432
rect 454866 627332 454990 627432
rect 455090 627332 455214 627432
rect 455314 627332 455438 627432
rect 455538 627332 455662 627432
rect 455762 627332 455886 627432
rect 455986 627332 456010 627432
rect 449350 627208 456010 627332
rect 449350 627108 449390 627208
rect 449490 627108 449614 627208
rect 449714 627108 449838 627208
rect 449938 627108 450062 627208
rect 450162 627108 450286 627208
rect 450386 627108 450510 627208
rect 450610 627108 450734 627208
rect 450834 627108 450958 627208
rect 451058 627108 451182 627208
rect 451282 627108 451406 627208
rect 451506 627108 451630 627208
rect 451730 627108 451854 627208
rect 451954 627108 452078 627208
rect 452178 627108 452302 627208
rect 452402 627108 452526 627208
rect 452626 627108 452750 627208
rect 452850 627108 452974 627208
rect 453074 627108 453198 627208
rect 453298 627108 453422 627208
rect 453522 627108 453646 627208
rect 453746 627108 453870 627208
rect 453970 627108 454094 627208
rect 454194 627108 454318 627208
rect 454418 627108 454542 627208
rect 454642 627108 454766 627208
rect 454866 627108 454990 627208
rect 455090 627108 455214 627208
rect 455314 627108 455438 627208
rect 455538 627108 455662 627208
rect 455762 627108 455886 627208
rect 455986 627108 456010 627208
rect 449350 626984 456010 627108
rect 449350 626884 449390 626984
rect 449490 626884 449614 626984
rect 449714 626884 449838 626984
rect 449938 626884 450062 626984
rect 450162 626884 450286 626984
rect 450386 626884 450510 626984
rect 450610 626884 450734 626984
rect 450834 626884 450958 626984
rect 451058 626884 451182 626984
rect 451282 626884 451406 626984
rect 451506 626884 451630 626984
rect 451730 626884 451854 626984
rect 451954 626884 452078 626984
rect 452178 626884 452302 626984
rect 452402 626884 452526 626984
rect 452626 626884 452750 626984
rect 452850 626884 452974 626984
rect 453074 626884 453198 626984
rect 453298 626884 453422 626984
rect 453522 626884 453646 626984
rect 453746 626884 453870 626984
rect 453970 626884 454094 626984
rect 454194 626884 454318 626984
rect 454418 626884 454542 626984
rect 454642 626884 454766 626984
rect 454866 626884 454990 626984
rect 455090 626884 455214 626984
rect 455314 626884 455438 626984
rect 455538 626884 455662 626984
rect 455762 626884 455886 626984
rect 455986 626884 456010 626984
rect 449350 626760 456010 626884
rect 449350 626660 449390 626760
rect 449490 626660 449614 626760
rect 449714 626660 449838 626760
rect 449938 626660 450062 626760
rect 450162 626660 450286 626760
rect 450386 626660 450510 626760
rect 450610 626660 450734 626760
rect 450834 626660 450958 626760
rect 451058 626660 451182 626760
rect 451282 626660 451406 626760
rect 451506 626660 451630 626760
rect 451730 626660 451854 626760
rect 451954 626660 452078 626760
rect 452178 626660 452302 626760
rect 452402 626660 452526 626760
rect 452626 626660 452750 626760
rect 452850 626660 452974 626760
rect 453074 626660 453198 626760
rect 453298 626660 453422 626760
rect 453522 626660 453646 626760
rect 453746 626660 453870 626760
rect 453970 626660 454094 626760
rect 454194 626660 454318 626760
rect 454418 626660 454542 626760
rect 454642 626660 454766 626760
rect 454866 626660 454990 626760
rect 455090 626660 455214 626760
rect 455314 626660 455438 626760
rect 455538 626660 455662 626760
rect 455762 626660 455886 626760
rect 455986 626660 456010 626760
rect 449350 626626 456010 626660
rect 475620 627676 482280 627706
rect 475620 627576 475660 627676
rect 475760 627576 475884 627676
rect 475984 627576 476108 627676
rect 476208 627576 476332 627676
rect 476432 627576 476556 627676
rect 476656 627576 476780 627676
rect 476880 627576 477004 627676
rect 477104 627576 477228 627676
rect 477328 627576 477452 627676
rect 477552 627576 477676 627676
rect 477776 627576 477900 627676
rect 478000 627576 478124 627676
rect 478224 627576 478348 627676
rect 478448 627576 478572 627676
rect 478672 627576 478796 627676
rect 478896 627576 479020 627676
rect 479120 627576 479244 627676
rect 479344 627576 479468 627676
rect 479568 627576 479692 627676
rect 479792 627576 479916 627676
rect 480016 627576 480140 627676
rect 480240 627576 480364 627676
rect 480464 627576 480588 627676
rect 480688 627576 480812 627676
rect 480912 627576 481036 627676
rect 481136 627576 481260 627676
rect 481360 627576 481484 627676
rect 481584 627576 481708 627676
rect 481808 627576 481932 627676
rect 482032 627576 482156 627676
rect 482256 627576 482280 627676
rect 475620 627452 482280 627576
rect 475620 627352 475660 627452
rect 475760 627352 475884 627452
rect 475984 627352 476108 627452
rect 476208 627352 476332 627452
rect 476432 627352 476556 627452
rect 476656 627352 476780 627452
rect 476880 627352 477004 627452
rect 477104 627352 477228 627452
rect 477328 627352 477452 627452
rect 477552 627352 477676 627452
rect 477776 627352 477900 627452
rect 478000 627352 478124 627452
rect 478224 627352 478348 627452
rect 478448 627352 478572 627452
rect 478672 627352 478796 627452
rect 478896 627352 479020 627452
rect 479120 627352 479244 627452
rect 479344 627352 479468 627452
rect 479568 627352 479692 627452
rect 479792 627352 479916 627452
rect 480016 627352 480140 627452
rect 480240 627352 480364 627452
rect 480464 627352 480588 627452
rect 480688 627352 480812 627452
rect 480912 627352 481036 627452
rect 481136 627352 481260 627452
rect 481360 627352 481484 627452
rect 481584 627352 481708 627452
rect 481808 627352 481932 627452
rect 482032 627352 482156 627452
rect 482256 627352 482280 627452
rect 475620 627228 482280 627352
rect 475620 627128 475660 627228
rect 475760 627128 475884 627228
rect 475984 627128 476108 627228
rect 476208 627128 476332 627228
rect 476432 627128 476556 627228
rect 476656 627128 476780 627228
rect 476880 627128 477004 627228
rect 477104 627128 477228 627228
rect 477328 627128 477452 627228
rect 477552 627128 477676 627228
rect 477776 627128 477900 627228
rect 478000 627128 478124 627228
rect 478224 627128 478348 627228
rect 478448 627128 478572 627228
rect 478672 627128 478796 627228
rect 478896 627128 479020 627228
rect 479120 627128 479244 627228
rect 479344 627128 479468 627228
rect 479568 627128 479692 627228
rect 479792 627128 479916 627228
rect 480016 627128 480140 627228
rect 480240 627128 480364 627228
rect 480464 627128 480588 627228
rect 480688 627128 480812 627228
rect 480912 627128 481036 627228
rect 481136 627128 481260 627228
rect 481360 627128 481484 627228
rect 481584 627128 481708 627228
rect 481808 627128 481932 627228
rect 482032 627128 482156 627228
rect 482256 627128 482280 627228
rect 475620 627004 482280 627128
rect 475620 626904 475660 627004
rect 475760 626904 475884 627004
rect 475984 626904 476108 627004
rect 476208 626904 476332 627004
rect 476432 626904 476556 627004
rect 476656 626904 476780 627004
rect 476880 626904 477004 627004
rect 477104 626904 477228 627004
rect 477328 626904 477452 627004
rect 477552 626904 477676 627004
rect 477776 626904 477900 627004
rect 478000 626904 478124 627004
rect 478224 626904 478348 627004
rect 478448 626904 478572 627004
rect 478672 626904 478796 627004
rect 478896 626904 479020 627004
rect 479120 626904 479244 627004
rect 479344 626904 479468 627004
rect 479568 626904 479692 627004
rect 479792 626904 479916 627004
rect 480016 626904 480140 627004
rect 480240 626904 480364 627004
rect 480464 626904 480588 627004
rect 480688 626904 480812 627004
rect 480912 626904 481036 627004
rect 481136 626904 481260 627004
rect 481360 626904 481484 627004
rect 481584 626904 481708 627004
rect 481808 626904 481932 627004
rect 482032 626904 482156 627004
rect 482256 626904 482280 627004
rect 475620 626780 482280 626904
rect 475620 626680 475660 626780
rect 475760 626680 475884 626780
rect 475984 626680 476108 626780
rect 476208 626680 476332 626780
rect 476432 626680 476556 626780
rect 476656 626680 476780 626780
rect 476880 626680 477004 626780
rect 477104 626680 477228 626780
rect 477328 626680 477452 626780
rect 477552 626680 477676 626780
rect 477776 626680 477900 626780
rect 478000 626680 478124 626780
rect 478224 626680 478348 626780
rect 478448 626680 478572 626780
rect 478672 626680 478796 626780
rect 478896 626680 479020 626780
rect 479120 626680 479244 626780
rect 479344 626680 479468 626780
rect 479568 626680 479692 626780
rect 479792 626680 479916 626780
rect 480016 626680 480140 626780
rect 480240 626680 480364 626780
rect 480464 626680 480588 626780
rect 480688 626680 480812 626780
rect 480912 626680 481036 626780
rect 481136 626680 481260 626780
rect 481360 626680 481484 626780
rect 481584 626680 481708 626780
rect 481808 626680 481932 626780
rect 482032 626680 482156 626780
rect 482256 626680 482280 626780
rect 475620 626646 482280 626680
<< via2 >>
rect 438920 654776 439020 654876
rect 439144 654776 439244 654876
rect 439368 654776 439468 654876
rect 439592 654776 439692 654876
rect 439816 654776 439916 654876
rect 440040 654776 440140 654876
rect 440264 654776 440364 654876
rect 440488 654776 440588 654876
rect 440712 654776 440812 654876
rect 440936 654776 441036 654876
rect 441160 654776 441260 654876
rect 441384 654776 441484 654876
rect 441608 654776 441708 654876
rect 441832 654776 441932 654876
rect 442056 654776 442156 654876
rect 442280 654776 442380 654876
rect 442504 654776 442604 654876
rect 442728 654776 442828 654876
rect 442952 654776 443052 654876
rect 443176 654776 443276 654876
rect 443400 654776 443500 654876
rect 443624 654776 443724 654876
rect 443848 654776 443948 654876
rect 444072 654776 444172 654876
rect 444296 654776 444396 654876
rect 444520 654776 444620 654876
rect 444744 654776 444844 654876
rect 444968 654776 445068 654876
rect 445192 654776 445292 654876
rect 445416 654776 445516 654876
rect 438920 654552 439020 654652
rect 439144 654552 439244 654652
rect 439368 654552 439468 654652
rect 439592 654552 439692 654652
rect 439816 654552 439916 654652
rect 440040 654552 440140 654652
rect 440264 654552 440364 654652
rect 440488 654552 440588 654652
rect 440712 654552 440812 654652
rect 440936 654552 441036 654652
rect 441160 654552 441260 654652
rect 441384 654552 441484 654652
rect 441608 654552 441708 654652
rect 441832 654552 441932 654652
rect 442056 654552 442156 654652
rect 442280 654552 442380 654652
rect 442504 654552 442604 654652
rect 442728 654552 442828 654652
rect 442952 654552 443052 654652
rect 443176 654552 443276 654652
rect 443400 654552 443500 654652
rect 443624 654552 443724 654652
rect 443848 654552 443948 654652
rect 444072 654552 444172 654652
rect 444296 654552 444396 654652
rect 444520 654552 444620 654652
rect 444744 654552 444844 654652
rect 444968 654552 445068 654652
rect 445192 654552 445292 654652
rect 445416 654552 445516 654652
rect 438920 654328 439020 654428
rect 439144 654328 439244 654428
rect 439368 654328 439468 654428
rect 439592 654328 439692 654428
rect 439816 654328 439916 654428
rect 440040 654328 440140 654428
rect 440264 654328 440364 654428
rect 440488 654328 440588 654428
rect 440712 654328 440812 654428
rect 440936 654328 441036 654428
rect 441160 654328 441260 654428
rect 441384 654328 441484 654428
rect 441608 654328 441708 654428
rect 441832 654328 441932 654428
rect 442056 654328 442156 654428
rect 442280 654328 442380 654428
rect 442504 654328 442604 654428
rect 442728 654328 442828 654428
rect 442952 654328 443052 654428
rect 443176 654328 443276 654428
rect 443400 654328 443500 654428
rect 443624 654328 443724 654428
rect 443848 654328 443948 654428
rect 444072 654328 444172 654428
rect 444296 654328 444396 654428
rect 444520 654328 444620 654428
rect 444744 654328 444844 654428
rect 444968 654328 445068 654428
rect 445192 654328 445292 654428
rect 445416 654328 445516 654428
rect 438920 654104 439020 654204
rect 439144 654104 439244 654204
rect 439368 654104 439468 654204
rect 439592 654104 439692 654204
rect 439816 654104 439916 654204
rect 440040 654104 440140 654204
rect 440264 654104 440364 654204
rect 440488 654104 440588 654204
rect 440712 654104 440812 654204
rect 440936 654104 441036 654204
rect 441160 654104 441260 654204
rect 441384 654104 441484 654204
rect 441608 654104 441708 654204
rect 441832 654104 441932 654204
rect 442056 654104 442156 654204
rect 442280 654104 442380 654204
rect 442504 654104 442604 654204
rect 442728 654104 442828 654204
rect 442952 654104 443052 654204
rect 443176 654104 443276 654204
rect 443400 654104 443500 654204
rect 443624 654104 443724 654204
rect 443848 654104 443948 654204
rect 444072 654104 444172 654204
rect 444296 654104 444396 654204
rect 444520 654104 444620 654204
rect 444744 654104 444844 654204
rect 444968 654104 445068 654204
rect 445192 654104 445292 654204
rect 445416 654104 445516 654204
rect 438920 653880 439020 653980
rect 439144 653880 439244 653980
rect 439368 653880 439468 653980
rect 439592 653880 439692 653980
rect 439816 653880 439916 653980
rect 440040 653880 440140 653980
rect 440264 653880 440364 653980
rect 440488 653880 440588 653980
rect 440712 653880 440812 653980
rect 440936 653880 441036 653980
rect 441160 653880 441260 653980
rect 441384 653880 441484 653980
rect 441608 653880 441708 653980
rect 441832 653880 441932 653980
rect 442056 653880 442156 653980
rect 442280 653880 442380 653980
rect 442504 653880 442604 653980
rect 442728 653880 442828 653980
rect 442952 653880 443052 653980
rect 443176 653880 443276 653980
rect 443400 653880 443500 653980
rect 443624 653880 443724 653980
rect 443848 653880 443948 653980
rect 444072 653880 444172 653980
rect 444296 653880 444396 653980
rect 444520 653880 444620 653980
rect 444744 653880 444844 653980
rect 444968 653880 445068 653980
rect 445192 653880 445292 653980
rect 445416 653880 445516 653980
rect 449390 654776 449490 654876
rect 449614 654776 449714 654876
rect 449838 654776 449938 654876
rect 450062 654776 450162 654876
rect 450286 654776 450386 654876
rect 450510 654776 450610 654876
rect 450734 654776 450834 654876
rect 450958 654776 451058 654876
rect 451182 654776 451282 654876
rect 451406 654776 451506 654876
rect 451630 654776 451730 654876
rect 451854 654776 451954 654876
rect 452078 654776 452178 654876
rect 452302 654776 452402 654876
rect 452526 654776 452626 654876
rect 452750 654776 452850 654876
rect 452974 654776 453074 654876
rect 453198 654776 453298 654876
rect 453422 654776 453522 654876
rect 453646 654776 453746 654876
rect 453870 654776 453970 654876
rect 454094 654776 454194 654876
rect 454318 654776 454418 654876
rect 454542 654776 454642 654876
rect 454766 654776 454866 654876
rect 454990 654776 455090 654876
rect 455214 654776 455314 654876
rect 455438 654776 455538 654876
rect 455662 654776 455762 654876
rect 455886 654776 455986 654876
rect 449390 654552 449490 654652
rect 449614 654552 449714 654652
rect 449838 654552 449938 654652
rect 450062 654552 450162 654652
rect 450286 654552 450386 654652
rect 450510 654552 450610 654652
rect 450734 654552 450834 654652
rect 450958 654552 451058 654652
rect 451182 654552 451282 654652
rect 451406 654552 451506 654652
rect 451630 654552 451730 654652
rect 451854 654552 451954 654652
rect 452078 654552 452178 654652
rect 452302 654552 452402 654652
rect 452526 654552 452626 654652
rect 452750 654552 452850 654652
rect 452974 654552 453074 654652
rect 453198 654552 453298 654652
rect 453422 654552 453522 654652
rect 453646 654552 453746 654652
rect 453870 654552 453970 654652
rect 454094 654552 454194 654652
rect 454318 654552 454418 654652
rect 454542 654552 454642 654652
rect 454766 654552 454866 654652
rect 454990 654552 455090 654652
rect 455214 654552 455314 654652
rect 455438 654552 455538 654652
rect 455662 654552 455762 654652
rect 455886 654552 455986 654652
rect 449390 654328 449490 654428
rect 449614 654328 449714 654428
rect 449838 654328 449938 654428
rect 450062 654328 450162 654428
rect 450286 654328 450386 654428
rect 450510 654328 450610 654428
rect 450734 654328 450834 654428
rect 450958 654328 451058 654428
rect 451182 654328 451282 654428
rect 451406 654328 451506 654428
rect 451630 654328 451730 654428
rect 451854 654328 451954 654428
rect 452078 654328 452178 654428
rect 452302 654328 452402 654428
rect 452526 654328 452626 654428
rect 452750 654328 452850 654428
rect 452974 654328 453074 654428
rect 453198 654328 453298 654428
rect 453422 654328 453522 654428
rect 453646 654328 453746 654428
rect 453870 654328 453970 654428
rect 454094 654328 454194 654428
rect 454318 654328 454418 654428
rect 454542 654328 454642 654428
rect 454766 654328 454866 654428
rect 454990 654328 455090 654428
rect 455214 654328 455314 654428
rect 455438 654328 455538 654428
rect 455662 654328 455762 654428
rect 455886 654328 455986 654428
rect 449390 654104 449490 654204
rect 449614 654104 449714 654204
rect 449838 654104 449938 654204
rect 450062 654104 450162 654204
rect 450286 654104 450386 654204
rect 450510 654104 450610 654204
rect 450734 654104 450834 654204
rect 450958 654104 451058 654204
rect 451182 654104 451282 654204
rect 451406 654104 451506 654204
rect 451630 654104 451730 654204
rect 451854 654104 451954 654204
rect 452078 654104 452178 654204
rect 452302 654104 452402 654204
rect 452526 654104 452626 654204
rect 452750 654104 452850 654204
rect 452974 654104 453074 654204
rect 453198 654104 453298 654204
rect 453422 654104 453522 654204
rect 453646 654104 453746 654204
rect 453870 654104 453970 654204
rect 454094 654104 454194 654204
rect 454318 654104 454418 654204
rect 454542 654104 454642 654204
rect 454766 654104 454866 654204
rect 454990 654104 455090 654204
rect 455214 654104 455314 654204
rect 455438 654104 455538 654204
rect 455662 654104 455762 654204
rect 455886 654104 455986 654204
rect 449390 653880 449490 653980
rect 449614 653880 449714 653980
rect 449838 653880 449938 653980
rect 450062 653880 450162 653980
rect 450286 653880 450386 653980
rect 450510 653880 450610 653980
rect 450734 653880 450834 653980
rect 450958 653880 451058 653980
rect 451182 653880 451282 653980
rect 451406 653880 451506 653980
rect 451630 653880 451730 653980
rect 451854 653880 451954 653980
rect 452078 653880 452178 653980
rect 452302 653880 452402 653980
rect 452526 653880 452626 653980
rect 452750 653880 452850 653980
rect 452974 653880 453074 653980
rect 453198 653880 453298 653980
rect 453422 653880 453522 653980
rect 453646 653880 453746 653980
rect 453870 653880 453970 653980
rect 454094 653880 454194 653980
rect 454318 653880 454418 653980
rect 454542 653880 454642 653980
rect 454766 653880 454866 653980
rect 454990 653880 455090 653980
rect 455214 653880 455314 653980
rect 455438 653880 455538 653980
rect 455662 653880 455762 653980
rect 455886 653880 455986 653980
rect 475660 654796 475760 654896
rect 475884 654796 475984 654896
rect 476108 654796 476208 654896
rect 476332 654796 476432 654896
rect 476556 654796 476656 654896
rect 476780 654796 476880 654896
rect 477004 654796 477104 654896
rect 477228 654796 477328 654896
rect 477452 654796 477552 654896
rect 477676 654796 477776 654896
rect 477900 654796 478000 654896
rect 478124 654796 478224 654896
rect 478348 654796 478448 654896
rect 478572 654796 478672 654896
rect 478796 654796 478896 654896
rect 479020 654796 479120 654896
rect 479244 654796 479344 654896
rect 479468 654796 479568 654896
rect 479692 654796 479792 654896
rect 479916 654796 480016 654896
rect 480140 654796 480240 654896
rect 480364 654796 480464 654896
rect 480588 654796 480688 654896
rect 480812 654796 480912 654896
rect 481036 654796 481136 654896
rect 481260 654796 481360 654896
rect 481484 654796 481584 654896
rect 481708 654796 481808 654896
rect 481932 654796 482032 654896
rect 482156 654796 482256 654896
rect 475660 654572 475760 654672
rect 475884 654572 475984 654672
rect 476108 654572 476208 654672
rect 476332 654572 476432 654672
rect 476556 654572 476656 654672
rect 476780 654572 476880 654672
rect 477004 654572 477104 654672
rect 477228 654572 477328 654672
rect 477452 654572 477552 654672
rect 477676 654572 477776 654672
rect 477900 654572 478000 654672
rect 478124 654572 478224 654672
rect 478348 654572 478448 654672
rect 478572 654572 478672 654672
rect 478796 654572 478896 654672
rect 479020 654572 479120 654672
rect 479244 654572 479344 654672
rect 479468 654572 479568 654672
rect 479692 654572 479792 654672
rect 479916 654572 480016 654672
rect 480140 654572 480240 654672
rect 480364 654572 480464 654672
rect 480588 654572 480688 654672
rect 480812 654572 480912 654672
rect 481036 654572 481136 654672
rect 481260 654572 481360 654672
rect 481484 654572 481584 654672
rect 481708 654572 481808 654672
rect 481932 654572 482032 654672
rect 482156 654572 482256 654672
rect 475660 654348 475760 654448
rect 475884 654348 475984 654448
rect 476108 654348 476208 654448
rect 476332 654348 476432 654448
rect 476556 654348 476656 654448
rect 476780 654348 476880 654448
rect 477004 654348 477104 654448
rect 477228 654348 477328 654448
rect 477452 654348 477552 654448
rect 477676 654348 477776 654448
rect 477900 654348 478000 654448
rect 478124 654348 478224 654448
rect 478348 654348 478448 654448
rect 478572 654348 478672 654448
rect 478796 654348 478896 654448
rect 479020 654348 479120 654448
rect 479244 654348 479344 654448
rect 479468 654348 479568 654448
rect 479692 654348 479792 654448
rect 479916 654348 480016 654448
rect 480140 654348 480240 654448
rect 480364 654348 480464 654448
rect 480588 654348 480688 654448
rect 480812 654348 480912 654448
rect 481036 654348 481136 654448
rect 481260 654348 481360 654448
rect 481484 654348 481584 654448
rect 481708 654348 481808 654448
rect 481932 654348 482032 654448
rect 482156 654348 482256 654448
rect 475660 654124 475760 654224
rect 475884 654124 475984 654224
rect 476108 654124 476208 654224
rect 476332 654124 476432 654224
rect 476556 654124 476656 654224
rect 476780 654124 476880 654224
rect 477004 654124 477104 654224
rect 477228 654124 477328 654224
rect 477452 654124 477552 654224
rect 477676 654124 477776 654224
rect 477900 654124 478000 654224
rect 478124 654124 478224 654224
rect 478348 654124 478448 654224
rect 478572 654124 478672 654224
rect 478796 654124 478896 654224
rect 479020 654124 479120 654224
rect 479244 654124 479344 654224
rect 479468 654124 479568 654224
rect 479692 654124 479792 654224
rect 479916 654124 480016 654224
rect 480140 654124 480240 654224
rect 480364 654124 480464 654224
rect 480588 654124 480688 654224
rect 480812 654124 480912 654224
rect 481036 654124 481136 654224
rect 481260 654124 481360 654224
rect 481484 654124 481584 654224
rect 481708 654124 481808 654224
rect 481932 654124 482032 654224
rect 482156 654124 482256 654224
rect 475660 653900 475760 654000
rect 475884 653900 475984 654000
rect 476108 653900 476208 654000
rect 476332 653900 476432 654000
rect 476556 653900 476656 654000
rect 476780 653900 476880 654000
rect 477004 653900 477104 654000
rect 477228 653900 477328 654000
rect 477452 653900 477552 654000
rect 477676 653900 477776 654000
rect 477900 653900 478000 654000
rect 478124 653900 478224 654000
rect 478348 653900 478448 654000
rect 478572 653900 478672 654000
rect 478796 653900 478896 654000
rect 479020 653900 479120 654000
rect 479244 653900 479344 654000
rect 479468 653900 479568 654000
rect 479692 653900 479792 654000
rect 479916 653900 480016 654000
rect 480140 653900 480240 654000
rect 480364 653900 480464 654000
rect 480588 653900 480688 654000
rect 480812 653900 480912 654000
rect 481036 653900 481136 654000
rect 481260 653900 481360 654000
rect 481484 653900 481584 654000
rect 481708 653900 481808 654000
rect 481932 653900 482032 654000
rect 482156 653900 482256 654000
rect 440696 652754 451952 652760
rect 440696 651928 440702 652754
rect 440702 651928 451946 652754
rect 451946 651928 451952 652754
rect 440696 651922 451952 651928
rect 437894 650078 437994 650178
rect 438118 650078 438218 650178
rect 438342 650078 438442 650178
rect 438566 650078 438666 650178
rect 438790 650078 438890 650178
rect 437894 649854 437994 649954
rect 438118 649854 438218 649954
rect 438342 649854 438442 649954
rect 438566 649854 438666 649954
rect 438790 649854 438890 649954
rect 437894 649630 437994 649730
rect 438118 649630 438218 649730
rect 438342 649630 438442 649730
rect 438566 649630 438666 649730
rect 438790 649630 438890 649730
rect 437894 649406 437994 649506
rect 438118 649406 438218 649506
rect 438342 649406 438442 649506
rect 438566 649406 438666 649506
rect 438790 649406 438890 649506
rect 437894 649182 437994 649282
rect 438118 649182 438218 649282
rect 438342 649182 438442 649282
rect 438566 649182 438666 649282
rect 438790 649182 438890 649282
rect 437894 648958 437994 649058
rect 438118 648958 438218 649058
rect 438342 648958 438442 649058
rect 438566 648958 438666 649058
rect 438790 648958 438890 649058
rect 437894 648734 437994 648834
rect 438118 648734 438218 648834
rect 438342 648734 438442 648834
rect 438566 648734 438666 648834
rect 438790 648734 438890 648834
rect 437894 648510 437994 648610
rect 438118 648510 438218 648610
rect 438342 648510 438442 648610
rect 438566 648510 438666 648610
rect 438790 648510 438890 648610
rect 437894 648286 437994 648386
rect 438118 648286 438218 648386
rect 438342 648286 438442 648386
rect 438566 648286 438666 648386
rect 438790 648286 438890 648386
rect 437894 648062 437994 648162
rect 438118 648062 438218 648162
rect 438342 648062 438442 648162
rect 438566 648062 438666 648162
rect 438790 648062 438890 648162
rect 437894 647838 437994 647938
rect 438118 647838 438218 647938
rect 438342 647838 438442 647938
rect 438566 647838 438666 647938
rect 438790 647838 438890 647938
rect 437894 647614 437994 647714
rect 438118 647614 438218 647714
rect 438342 647614 438442 647714
rect 438566 647614 438666 647714
rect 438790 647614 438890 647714
rect 437894 647390 437994 647490
rect 438118 647390 438218 647490
rect 438342 647390 438442 647490
rect 438566 647390 438666 647490
rect 438790 647390 438890 647490
rect 437894 647166 437994 647266
rect 438118 647166 438218 647266
rect 438342 647166 438442 647266
rect 438566 647166 438666 647266
rect 438790 647166 438890 647266
rect 437894 646942 437994 647042
rect 438118 646942 438218 647042
rect 438342 646942 438442 647042
rect 438566 646942 438666 647042
rect 438790 646942 438890 647042
rect 437894 646718 437994 646818
rect 438118 646718 438218 646818
rect 438342 646718 438442 646818
rect 438566 646718 438666 646818
rect 438790 646718 438890 646818
rect 437894 646494 437994 646594
rect 438118 646494 438218 646594
rect 438342 646494 438442 646594
rect 438566 646494 438666 646594
rect 438790 646494 438890 646594
rect 437894 646270 437994 646370
rect 438118 646270 438218 646370
rect 438342 646270 438442 646370
rect 438566 646270 438666 646370
rect 438790 646270 438890 646370
rect 482174 650078 482274 650178
rect 482398 650078 482498 650178
rect 482622 650078 482722 650178
rect 482846 650078 482946 650178
rect 483070 650078 483170 650178
rect 482174 649854 482274 649954
rect 482398 649854 482498 649954
rect 482622 649854 482722 649954
rect 482846 649854 482946 649954
rect 483070 649854 483170 649954
rect 482174 649630 482274 649730
rect 482398 649630 482498 649730
rect 482622 649630 482722 649730
rect 482846 649630 482946 649730
rect 483070 649630 483170 649730
rect 482174 649406 482274 649506
rect 482398 649406 482498 649506
rect 482622 649406 482722 649506
rect 482846 649406 482946 649506
rect 483070 649406 483170 649506
rect 482174 649182 482274 649282
rect 482398 649182 482498 649282
rect 482622 649182 482722 649282
rect 482846 649182 482946 649282
rect 483070 649182 483170 649282
rect 482174 648958 482274 649058
rect 482398 648958 482498 649058
rect 482622 648958 482722 649058
rect 482846 648958 482946 649058
rect 483070 648958 483170 649058
rect 482174 648734 482274 648834
rect 482398 648734 482498 648834
rect 482622 648734 482722 648834
rect 482846 648734 482946 648834
rect 483070 648734 483170 648834
rect 482174 648510 482274 648610
rect 482398 648510 482498 648610
rect 482622 648510 482722 648610
rect 482846 648510 482946 648610
rect 483070 648510 483170 648610
rect 482174 648286 482274 648386
rect 482398 648286 482498 648386
rect 482622 648286 482722 648386
rect 482846 648286 482946 648386
rect 483070 648286 483170 648386
rect 482174 648062 482274 648162
rect 482398 648062 482498 648162
rect 482622 648062 482722 648162
rect 482846 648062 482946 648162
rect 483070 648062 483170 648162
rect 482174 647838 482274 647938
rect 482398 647838 482498 647938
rect 482622 647838 482722 647938
rect 482846 647838 482946 647938
rect 483070 647838 483170 647938
rect 482174 647614 482274 647714
rect 482398 647614 482498 647714
rect 482622 647614 482722 647714
rect 482846 647614 482946 647714
rect 483070 647614 483170 647714
rect 482174 647390 482274 647490
rect 482398 647390 482498 647490
rect 482622 647390 482722 647490
rect 482846 647390 482946 647490
rect 483070 647390 483170 647490
rect 482174 647166 482274 647266
rect 482398 647166 482498 647266
rect 482622 647166 482722 647266
rect 482846 647166 482946 647266
rect 483070 647166 483170 647266
rect 482174 646942 482274 647042
rect 482398 646942 482498 647042
rect 482622 646942 482722 647042
rect 482846 646942 482946 647042
rect 483070 646942 483170 647042
rect 437894 646046 437994 646146
rect 438118 646046 438218 646146
rect 438342 646046 438442 646146
rect 438566 646046 438666 646146
rect 438790 646046 438890 646146
rect 437894 645822 437994 645922
rect 438118 645822 438218 645922
rect 438342 645822 438442 645922
rect 438566 645822 438666 645922
rect 438790 645822 438890 645922
rect 437894 645598 437994 645698
rect 438118 645598 438218 645698
rect 438342 645598 438442 645698
rect 438566 645598 438666 645698
rect 438790 645598 438890 645698
rect 437894 645374 437994 645474
rect 438118 645374 438218 645474
rect 438342 645374 438442 645474
rect 438566 645374 438666 645474
rect 438790 645374 438890 645474
rect 437894 645150 437994 645250
rect 438118 645150 438218 645250
rect 438342 645150 438442 645250
rect 438566 645150 438666 645250
rect 438790 645150 438890 645250
rect 437894 644926 437994 645026
rect 438118 644926 438218 645026
rect 438342 644926 438442 645026
rect 438566 644926 438666 645026
rect 438790 644926 438890 645026
rect 437894 644702 437994 644802
rect 438118 644702 438218 644802
rect 438342 644702 438442 644802
rect 438566 644702 438666 644802
rect 438790 644702 438890 644802
rect 437894 644478 437994 644578
rect 438118 644478 438218 644578
rect 438342 644478 438442 644578
rect 438566 644478 438666 644578
rect 438790 644478 438890 644578
rect 437894 644254 437994 644354
rect 438118 644254 438218 644354
rect 438342 644254 438442 644354
rect 438566 644254 438666 644354
rect 438790 644254 438890 644354
rect 437894 644030 437994 644130
rect 438118 644030 438218 644130
rect 438342 644030 438442 644130
rect 438566 644030 438666 644130
rect 438790 644030 438890 644130
rect 437894 643806 437994 643906
rect 438118 643806 438218 643906
rect 438342 643806 438442 643906
rect 438566 643806 438666 643906
rect 438790 643806 438890 643906
rect 437894 643582 437994 643682
rect 438118 643582 438218 643682
rect 438342 643582 438442 643682
rect 438566 643582 438666 643682
rect 438790 643582 438890 643682
rect 482174 646718 482274 646818
rect 482398 646718 482498 646818
rect 482622 646718 482722 646818
rect 482846 646718 482946 646818
rect 483070 646718 483170 646818
rect 482174 646494 482274 646594
rect 482398 646494 482498 646594
rect 482622 646494 482722 646594
rect 482846 646494 482946 646594
rect 483070 646494 483170 646594
rect 482174 646270 482274 646370
rect 482398 646270 482498 646370
rect 482622 646270 482722 646370
rect 482846 646270 482946 646370
rect 483070 646270 483170 646370
rect 482174 646046 482274 646146
rect 482398 646046 482498 646146
rect 482622 646046 482722 646146
rect 482846 646046 482946 646146
rect 483070 646046 483170 646146
rect 482174 645822 482274 645922
rect 482398 645822 482498 645922
rect 482622 645822 482722 645922
rect 482846 645822 482946 645922
rect 483070 645822 483170 645922
rect 482174 645598 482274 645698
rect 482398 645598 482498 645698
rect 482622 645598 482722 645698
rect 482846 645598 482946 645698
rect 483070 645598 483170 645698
rect 482174 645374 482274 645474
rect 482398 645374 482498 645474
rect 482622 645374 482722 645474
rect 482846 645374 482946 645474
rect 483070 645374 483170 645474
rect 482174 645150 482274 645250
rect 482398 645150 482498 645250
rect 482622 645150 482722 645250
rect 482846 645150 482946 645250
rect 483070 645150 483170 645250
rect 482174 644926 482274 645026
rect 482398 644926 482498 645026
rect 482622 644926 482722 645026
rect 482846 644926 482946 645026
rect 483070 644926 483170 645026
rect 482174 644702 482274 644802
rect 482398 644702 482498 644802
rect 482622 644702 482722 644802
rect 482846 644702 482946 644802
rect 483070 644702 483170 644802
rect 482174 644478 482274 644578
rect 482398 644478 482498 644578
rect 482622 644478 482722 644578
rect 482846 644478 482946 644578
rect 483070 644478 483170 644578
rect 482174 644254 482274 644354
rect 482398 644254 482498 644354
rect 482622 644254 482722 644354
rect 482846 644254 482946 644354
rect 483070 644254 483170 644354
rect 482174 644030 482274 644130
rect 482398 644030 482498 644130
rect 482622 644030 482722 644130
rect 482846 644030 482946 644130
rect 483070 644030 483170 644130
rect 482174 643806 482274 643906
rect 482398 643806 482498 643906
rect 482622 643806 482722 643906
rect 482846 643806 482946 643906
rect 483070 643806 483170 643906
rect 482174 643582 482274 643682
rect 482398 643582 482498 643682
rect 482622 643582 482722 643682
rect 482846 643582 482946 643682
rect 483070 643582 483170 643682
rect 459444 640850 459644 641050
rect 459878 640850 460078 641050
rect 460312 640850 460512 641050
rect 460746 640850 460946 641050
rect 461180 640850 461380 641050
rect 461614 640850 461814 641050
rect 462048 640850 462248 641050
rect 462482 640850 462682 641050
rect 462916 640850 463116 641050
rect 463350 640850 463550 641050
rect 463784 640850 463984 641050
rect 464184 640850 464384 641050
rect 464584 640850 464784 641050
rect 464984 640850 465184 641050
rect 465384 640850 465584 641050
rect 465784 640850 465984 641050
rect 466184 640850 466384 641050
rect 466584 640850 466784 641050
rect 466984 640850 467184 641050
rect 467384 640850 467584 641050
rect 459444 640416 459644 640616
rect 459878 640416 460078 640616
rect 460312 640416 460512 640616
rect 460746 640416 460946 640616
rect 461180 640416 461380 640616
rect 461614 640416 461814 640616
rect 462048 640416 462248 640616
rect 462482 640416 462682 640616
rect 462916 640416 463116 640616
rect 463350 640416 463550 640616
rect 463784 640416 463984 640616
rect 468984 640850 469184 641050
rect 469384 640850 469584 641050
rect 469784 640850 469984 641050
rect 470184 640850 470384 641050
rect 470584 640850 470784 641050
rect 470984 640850 471184 641050
rect 471384 640850 471584 641050
rect 471784 640850 471984 641050
rect 472184 640850 472384 641050
rect 459444 639982 459644 640182
rect 459878 639982 460078 640182
rect 460312 639982 460512 640182
rect 460746 639982 460946 640182
rect 461180 639982 461380 640182
rect 461614 639982 461814 640182
rect 462048 639982 462248 640182
rect 462482 639982 462682 640182
rect 462916 639982 463116 640182
rect 463350 639982 463550 640182
rect 463784 639982 463984 640182
rect 452996 639098 453864 639474
rect 453864 639098 455852 639474
rect 455852 639098 467564 639474
rect 467564 639098 469552 639474
rect 469552 639098 472876 639474
rect 472876 639098 473318 639474
rect 452996 638684 473318 639098
rect 452996 638490 453864 638684
rect 453864 638490 455852 638684
rect 455852 638490 467564 638684
rect 467564 638490 469552 638684
rect 469552 638490 473318 638684
rect 443024 638152 443084 638212
rect 443144 638152 443204 638212
rect 443264 638152 443324 638212
rect 443384 638152 443444 638212
rect 443504 638152 443564 638212
rect 443024 638032 443084 638092
rect 443144 638032 443204 638092
rect 443264 638032 443324 638092
rect 443384 638032 443444 638092
rect 443504 638032 443564 638092
rect 437894 636678 437994 636778
rect 438118 636678 438218 636778
rect 438342 636678 438442 636778
rect 438566 636678 438666 636778
rect 438790 636678 438890 636778
rect 437894 636454 437994 636554
rect 438118 636454 438218 636554
rect 438342 636454 438442 636554
rect 438566 636454 438666 636554
rect 438790 636454 438890 636554
rect 437894 636230 437994 636330
rect 438118 636230 438218 636330
rect 438342 636230 438442 636330
rect 438566 636230 438666 636330
rect 438790 636230 438890 636330
rect 482174 636678 482274 636778
rect 482398 636678 482498 636778
rect 482622 636678 482722 636778
rect 482846 636678 482946 636778
rect 483070 636678 483170 636778
rect 482174 636454 482274 636554
rect 482398 636454 482498 636554
rect 482622 636454 482722 636554
rect 482846 636454 482946 636554
rect 483070 636454 483170 636554
rect 482174 636230 482274 636330
rect 482398 636230 482498 636330
rect 482622 636230 482722 636330
rect 482846 636230 482946 636330
rect 483070 636230 483170 636330
rect 437894 636006 437994 636106
rect 438118 636006 438218 636106
rect 438342 636006 438442 636106
rect 438566 636006 438666 636106
rect 438790 636006 438890 636106
rect 437894 635782 437994 635882
rect 438118 635782 438218 635882
rect 438342 635782 438442 635882
rect 438566 635782 438666 635882
rect 438790 635782 438890 635882
rect 482174 636006 482274 636106
rect 482398 636006 482498 636106
rect 482622 636006 482722 636106
rect 482846 636006 482946 636106
rect 483070 636006 483170 636106
rect 482174 635782 482274 635882
rect 482398 635782 482498 635882
rect 482622 635782 482722 635882
rect 482846 635782 482946 635882
rect 483070 635782 483170 635882
rect 437894 635558 437994 635658
rect 438118 635558 438218 635658
rect 438342 635558 438442 635658
rect 438566 635558 438666 635658
rect 438790 635558 438890 635658
rect 437894 635334 437994 635434
rect 438118 635334 438218 635434
rect 438342 635334 438442 635434
rect 438566 635334 438666 635434
rect 438790 635334 438890 635434
rect 437894 635110 437994 635210
rect 438118 635110 438218 635210
rect 438342 635110 438442 635210
rect 438566 635110 438666 635210
rect 438790 635110 438890 635210
rect 482174 635558 482274 635658
rect 482398 635558 482498 635658
rect 482622 635558 482722 635658
rect 482846 635558 482946 635658
rect 483070 635558 483170 635658
rect 482174 635334 482274 635434
rect 482398 635334 482498 635434
rect 482622 635334 482722 635434
rect 482846 635334 482946 635434
rect 483070 635334 483170 635434
rect 482174 635110 482274 635210
rect 482398 635110 482498 635210
rect 482622 635110 482722 635210
rect 482846 635110 482946 635210
rect 483070 635110 483170 635210
rect 437894 634886 437994 634986
rect 438118 634886 438218 634986
rect 438342 634886 438442 634986
rect 438566 634886 438666 634986
rect 438790 634886 438890 634986
rect 437894 634662 437994 634762
rect 438118 634662 438218 634762
rect 438342 634662 438442 634762
rect 438566 634662 438666 634762
rect 438790 634662 438890 634762
rect 482174 634886 482274 634986
rect 482398 634886 482498 634986
rect 482622 634886 482722 634986
rect 482846 634886 482946 634986
rect 483070 634886 483170 634986
rect 482174 634662 482274 634762
rect 482398 634662 482498 634762
rect 482622 634662 482722 634762
rect 482846 634662 482946 634762
rect 483070 634662 483170 634762
rect 437894 634438 437994 634538
rect 438118 634438 438218 634538
rect 438342 634438 438442 634538
rect 438566 634438 438666 634538
rect 438790 634438 438890 634538
rect 437894 634214 437994 634314
rect 438118 634214 438218 634314
rect 438342 634214 438442 634314
rect 438566 634214 438666 634314
rect 438790 634214 438890 634314
rect 437894 633990 437994 634090
rect 438118 633990 438218 634090
rect 438342 633990 438442 634090
rect 438566 633990 438666 634090
rect 438790 633990 438890 634090
rect 437894 633766 437994 633866
rect 438118 633766 438218 633866
rect 438342 633766 438442 633866
rect 438566 633766 438666 633866
rect 438790 633766 438890 633866
rect 437894 633542 437994 633642
rect 438118 633542 438218 633642
rect 438342 633542 438442 633642
rect 438566 633542 438666 633642
rect 438790 633542 438890 633642
rect 437894 633318 437994 633418
rect 438118 633318 438218 633418
rect 438342 633318 438442 633418
rect 438566 633318 438666 633418
rect 438790 633318 438890 633418
rect 437894 633094 437994 633194
rect 438118 633094 438218 633194
rect 438342 633094 438442 633194
rect 438566 633094 438666 633194
rect 438790 633094 438890 633194
rect 437894 632870 437994 632970
rect 438118 632870 438218 632970
rect 438342 632870 438442 632970
rect 438566 632870 438666 632970
rect 438790 632870 438890 632970
rect 437894 632646 437994 632746
rect 438118 632646 438218 632746
rect 438342 632646 438442 632746
rect 438566 632646 438666 632746
rect 438790 632646 438890 632746
rect 482174 634438 482274 634538
rect 482398 634438 482498 634538
rect 482622 634438 482722 634538
rect 482846 634438 482946 634538
rect 483070 634438 483170 634538
rect 482174 634214 482274 634314
rect 482398 634214 482498 634314
rect 482622 634214 482722 634314
rect 482846 634214 482946 634314
rect 483070 634214 483170 634314
rect 482174 633990 482274 634090
rect 482398 633990 482498 634090
rect 482622 633990 482722 634090
rect 482846 633990 482946 634090
rect 483070 633990 483170 634090
rect 482174 633766 482274 633866
rect 482398 633766 482498 633866
rect 482622 633766 482722 633866
rect 482846 633766 482946 633866
rect 483070 633766 483170 633866
rect 482174 633542 482274 633642
rect 482398 633542 482498 633642
rect 482622 633542 482722 633642
rect 482846 633542 482946 633642
rect 483070 633542 483170 633642
rect 482174 633318 482274 633418
rect 482398 633318 482498 633418
rect 482622 633318 482722 633418
rect 482846 633318 482946 633418
rect 483070 633318 483170 633418
rect 482174 633094 482274 633194
rect 482398 633094 482498 633194
rect 482622 633094 482722 633194
rect 482846 633094 482946 633194
rect 483070 633094 483170 633194
rect 482174 632870 482274 632970
rect 482398 632870 482498 632970
rect 482622 632870 482722 632970
rect 482846 632870 482946 632970
rect 483070 632870 483170 632970
rect 482174 632646 482274 632746
rect 482398 632646 482498 632746
rect 482622 632646 482722 632746
rect 482846 632646 482946 632746
rect 483070 632646 483170 632746
rect 437894 632422 437994 632522
rect 438118 632422 438218 632522
rect 438342 632422 438442 632522
rect 438566 632422 438666 632522
rect 438790 632422 438890 632522
rect 482174 632422 482274 632522
rect 482398 632422 482498 632522
rect 482622 632422 482722 632522
rect 482846 632422 482946 632522
rect 483070 632422 483170 632522
rect 437894 632198 437994 632298
rect 438118 632198 438218 632298
rect 438342 632198 438442 632298
rect 438566 632198 438666 632298
rect 438790 632198 438890 632298
rect 437894 631974 437994 632074
rect 438118 631974 438218 632074
rect 438342 631974 438442 632074
rect 438566 631974 438666 632074
rect 438790 631974 438890 632074
rect 443648 632065 444248 632317
rect 452139 632065 452739 632317
rect 482174 632198 482274 632298
rect 482398 632198 482498 632298
rect 482622 632198 482722 632298
rect 482846 632198 482946 632298
rect 483070 632198 483170 632298
rect 482174 631974 482274 632074
rect 482398 631974 482498 632074
rect 482622 631974 482722 632074
rect 482846 631974 482946 632074
rect 483070 631974 483170 632074
rect 437894 631750 437994 631850
rect 438118 631750 438218 631850
rect 438342 631750 438442 631850
rect 438566 631750 438666 631850
rect 438790 631750 438890 631850
rect 437894 631526 437994 631626
rect 438118 631526 438218 631626
rect 438342 631526 438442 631626
rect 438566 631526 438666 631626
rect 438790 631526 438890 631626
rect 437894 631302 437994 631402
rect 438118 631302 438218 631402
rect 438342 631302 438442 631402
rect 438566 631302 438666 631402
rect 438790 631302 438890 631402
rect 437894 631078 437994 631178
rect 438118 631078 438218 631178
rect 438342 631078 438442 631178
rect 438566 631078 438666 631178
rect 438790 631078 438890 631178
rect 437894 630854 437994 630954
rect 438118 630854 438218 630954
rect 438342 630854 438442 630954
rect 438566 630854 438666 630954
rect 438790 630854 438890 630954
rect 482174 631750 482274 631850
rect 482398 631750 482498 631850
rect 482622 631750 482722 631850
rect 482846 631750 482946 631850
rect 483070 631750 483170 631850
rect 482174 631526 482274 631626
rect 482398 631526 482498 631626
rect 482622 631526 482722 631626
rect 482846 631526 482946 631626
rect 483070 631526 483170 631626
rect 482174 631302 482274 631402
rect 482398 631302 482498 631402
rect 482622 631302 482722 631402
rect 482846 631302 482946 631402
rect 483070 631302 483170 631402
rect 482174 631078 482274 631178
rect 482398 631078 482498 631178
rect 482622 631078 482722 631178
rect 482846 631078 482946 631178
rect 483070 631078 483170 631178
rect 437894 630630 437994 630730
rect 438118 630630 438218 630730
rect 438342 630630 438442 630730
rect 438566 630630 438666 630730
rect 438790 630630 438890 630730
rect 437894 630406 437994 630506
rect 438118 630406 438218 630506
rect 438342 630406 438442 630506
rect 438566 630406 438666 630506
rect 438790 630406 438890 630506
rect 437894 630182 437994 630282
rect 438118 630182 438218 630282
rect 438342 630182 438442 630282
rect 438566 630182 438666 630282
rect 438790 630182 438890 630282
rect 482174 630854 482274 630954
rect 482398 630854 482498 630954
rect 482622 630854 482722 630954
rect 482846 630854 482946 630954
rect 483070 630854 483170 630954
rect 482174 630630 482274 630730
rect 482398 630630 482498 630730
rect 482622 630630 482722 630730
rect 482846 630630 482946 630730
rect 483070 630630 483170 630730
rect 482174 630406 482274 630506
rect 482398 630406 482498 630506
rect 482622 630406 482722 630506
rect 482846 630406 482946 630506
rect 483070 630406 483170 630506
rect 482174 630182 482274 630282
rect 482398 630182 482498 630282
rect 482622 630182 482722 630282
rect 482846 630182 482946 630282
rect 483070 630182 483170 630282
rect 442990 629240 452236 629244
rect 442990 629136 443008 629240
rect 443008 629136 443060 629240
rect 443060 629136 443630 629240
rect 443630 629136 443682 629240
rect 443682 629136 444088 629240
rect 444088 629136 444140 629240
rect 444140 629136 444664 629240
rect 444664 629136 444716 629240
rect 444716 629136 445236 629240
rect 445236 629136 445288 629240
rect 445288 629136 445808 629240
rect 445808 629136 445860 629240
rect 445860 629136 446380 629240
rect 446380 629136 446432 629240
rect 446432 629136 446952 629240
rect 446952 629136 447004 629240
rect 447004 629136 447524 629240
rect 447524 629136 447576 629240
rect 447576 629136 448096 629240
rect 448096 629136 448148 629240
rect 448148 629136 448668 629240
rect 448668 629136 448720 629240
rect 448720 629136 449240 629240
rect 449240 629136 449292 629240
rect 449292 629136 449812 629240
rect 449812 629136 449864 629240
rect 449864 629136 450384 629240
rect 450384 629136 450436 629240
rect 450436 629136 450956 629240
rect 450956 629136 451008 629240
rect 451008 629136 451066 629240
rect 451066 629136 451118 629240
rect 451118 629136 451524 629240
rect 451524 629136 451576 629240
rect 451576 629136 452136 629240
rect 452136 629136 452188 629240
rect 452188 629136 452236 629240
rect 442990 629130 452236 629136
rect 452754 629010 470692 629012
rect 452754 628930 454338 629010
rect 454338 628930 454418 629010
rect 454418 628930 455258 629010
rect 455258 628930 455338 629010
rect 455338 628930 456178 629010
rect 456178 628930 456258 629010
rect 456258 628930 457098 629010
rect 457098 628930 457178 629010
rect 457178 628930 458018 629010
rect 458018 628930 458098 629010
rect 458098 628930 459838 629010
rect 459838 628930 459918 629010
rect 459918 628930 460758 629010
rect 460758 628930 460838 629010
rect 460838 628930 461678 629010
rect 461678 628930 461758 629010
rect 461758 628930 462598 629010
rect 462598 628930 462678 629010
rect 462678 628930 463518 629010
rect 463518 628930 463598 629010
rect 463598 628930 465338 629010
rect 465338 628930 465418 629010
rect 465418 628930 466258 629010
rect 466258 628930 466338 629010
rect 466338 628930 467178 629010
rect 467178 628930 467258 629010
rect 467258 628930 468098 629010
rect 468098 628930 468178 629010
rect 468178 628930 469018 629010
rect 469018 628930 469098 629010
rect 469098 628930 470692 629010
rect 452754 628890 470692 628930
rect 452754 628790 452848 628890
rect 452848 628790 453248 628890
rect 453248 628790 458758 628890
rect 458758 628790 459158 628890
rect 459158 628790 464258 628890
rect 464258 628790 464658 628890
rect 464658 628888 470692 628890
rect 464658 628790 470214 628888
rect 452754 628788 470214 628790
rect 470214 628788 470614 628888
rect 470614 628788 470692 628888
rect 452754 628694 470692 628788
rect 438920 627556 439020 627656
rect 439144 627556 439244 627656
rect 439368 627556 439468 627656
rect 439592 627556 439692 627656
rect 439816 627556 439916 627656
rect 440040 627556 440140 627656
rect 440264 627556 440364 627656
rect 440488 627556 440588 627656
rect 440712 627556 440812 627656
rect 440936 627556 441036 627656
rect 441160 627556 441260 627656
rect 441384 627556 441484 627656
rect 441608 627556 441708 627656
rect 441832 627556 441932 627656
rect 442056 627556 442156 627656
rect 442280 627556 442380 627656
rect 442504 627556 442604 627656
rect 442728 627556 442828 627656
rect 442952 627556 443052 627656
rect 443176 627556 443276 627656
rect 443400 627556 443500 627656
rect 443624 627556 443724 627656
rect 443848 627556 443948 627656
rect 444072 627556 444172 627656
rect 444296 627556 444396 627656
rect 444520 627556 444620 627656
rect 444744 627556 444844 627656
rect 444968 627556 445068 627656
rect 445192 627556 445292 627656
rect 445416 627556 445516 627656
rect 438920 627332 439020 627432
rect 439144 627332 439244 627432
rect 439368 627332 439468 627432
rect 439592 627332 439692 627432
rect 439816 627332 439916 627432
rect 440040 627332 440140 627432
rect 440264 627332 440364 627432
rect 440488 627332 440588 627432
rect 440712 627332 440812 627432
rect 440936 627332 441036 627432
rect 441160 627332 441260 627432
rect 441384 627332 441484 627432
rect 441608 627332 441708 627432
rect 441832 627332 441932 627432
rect 442056 627332 442156 627432
rect 442280 627332 442380 627432
rect 442504 627332 442604 627432
rect 442728 627332 442828 627432
rect 442952 627332 443052 627432
rect 443176 627332 443276 627432
rect 443400 627332 443500 627432
rect 443624 627332 443724 627432
rect 443848 627332 443948 627432
rect 444072 627332 444172 627432
rect 444296 627332 444396 627432
rect 444520 627332 444620 627432
rect 444744 627332 444844 627432
rect 444968 627332 445068 627432
rect 445192 627332 445292 627432
rect 445416 627332 445516 627432
rect 438920 627108 439020 627208
rect 439144 627108 439244 627208
rect 439368 627108 439468 627208
rect 439592 627108 439692 627208
rect 439816 627108 439916 627208
rect 440040 627108 440140 627208
rect 440264 627108 440364 627208
rect 440488 627108 440588 627208
rect 440712 627108 440812 627208
rect 440936 627108 441036 627208
rect 441160 627108 441260 627208
rect 441384 627108 441484 627208
rect 441608 627108 441708 627208
rect 441832 627108 441932 627208
rect 442056 627108 442156 627208
rect 442280 627108 442380 627208
rect 442504 627108 442604 627208
rect 442728 627108 442828 627208
rect 442952 627108 443052 627208
rect 443176 627108 443276 627208
rect 443400 627108 443500 627208
rect 443624 627108 443724 627208
rect 443848 627108 443948 627208
rect 444072 627108 444172 627208
rect 444296 627108 444396 627208
rect 444520 627108 444620 627208
rect 444744 627108 444844 627208
rect 444968 627108 445068 627208
rect 445192 627108 445292 627208
rect 445416 627108 445516 627208
rect 438920 626884 439020 626984
rect 439144 626884 439244 626984
rect 439368 626884 439468 626984
rect 439592 626884 439692 626984
rect 439816 626884 439916 626984
rect 440040 626884 440140 626984
rect 440264 626884 440364 626984
rect 440488 626884 440588 626984
rect 440712 626884 440812 626984
rect 440936 626884 441036 626984
rect 441160 626884 441260 626984
rect 441384 626884 441484 626984
rect 441608 626884 441708 626984
rect 441832 626884 441932 626984
rect 442056 626884 442156 626984
rect 442280 626884 442380 626984
rect 442504 626884 442604 626984
rect 442728 626884 442828 626984
rect 442952 626884 443052 626984
rect 443176 626884 443276 626984
rect 443400 626884 443500 626984
rect 443624 626884 443724 626984
rect 443848 626884 443948 626984
rect 444072 626884 444172 626984
rect 444296 626884 444396 626984
rect 444520 626884 444620 626984
rect 444744 626884 444844 626984
rect 444968 626884 445068 626984
rect 445192 626884 445292 626984
rect 445416 626884 445516 626984
rect 438920 626660 439020 626760
rect 439144 626660 439244 626760
rect 439368 626660 439468 626760
rect 439592 626660 439692 626760
rect 439816 626660 439916 626760
rect 440040 626660 440140 626760
rect 440264 626660 440364 626760
rect 440488 626660 440588 626760
rect 440712 626660 440812 626760
rect 440936 626660 441036 626760
rect 441160 626660 441260 626760
rect 441384 626660 441484 626760
rect 441608 626660 441708 626760
rect 441832 626660 441932 626760
rect 442056 626660 442156 626760
rect 442280 626660 442380 626760
rect 442504 626660 442604 626760
rect 442728 626660 442828 626760
rect 442952 626660 443052 626760
rect 443176 626660 443276 626760
rect 443400 626660 443500 626760
rect 443624 626660 443724 626760
rect 443848 626660 443948 626760
rect 444072 626660 444172 626760
rect 444296 626660 444396 626760
rect 444520 626660 444620 626760
rect 444744 626660 444844 626760
rect 444968 626660 445068 626760
rect 445192 626660 445292 626760
rect 445416 626660 445516 626760
rect 449390 627556 449490 627656
rect 449614 627556 449714 627656
rect 449838 627556 449938 627656
rect 450062 627556 450162 627656
rect 450286 627556 450386 627656
rect 450510 627556 450610 627656
rect 450734 627556 450834 627656
rect 450958 627556 451058 627656
rect 451182 627556 451282 627656
rect 451406 627556 451506 627656
rect 451630 627556 451730 627656
rect 451854 627556 451954 627656
rect 452078 627556 452178 627656
rect 452302 627556 452402 627656
rect 452526 627556 452626 627656
rect 452750 627556 452850 627656
rect 452974 627556 453074 627656
rect 453198 627556 453298 627656
rect 453422 627556 453522 627656
rect 453646 627556 453746 627656
rect 453870 627556 453970 627656
rect 454094 627556 454194 627656
rect 454318 627556 454418 627656
rect 454542 627556 454642 627656
rect 454766 627556 454866 627656
rect 454990 627556 455090 627656
rect 455214 627556 455314 627656
rect 455438 627556 455538 627656
rect 455662 627556 455762 627656
rect 455886 627556 455986 627656
rect 449390 627332 449490 627432
rect 449614 627332 449714 627432
rect 449838 627332 449938 627432
rect 450062 627332 450162 627432
rect 450286 627332 450386 627432
rect 450510 627332 450610 627432
rect 450734 627332 450834 627432
rect 450958 627332 451058 627432
rect 451182 627332 451282 627432
rect 451406 627332 451506 627432
rect 451630 627332 451730 627432
rect 451854 627332 451954 627432
rect 452078 627332 452178 627432
rect 452302 627332 452402 627432
rect 452526 627332 452626 627432
rect 452750 627332 452850 627432
rect 452974 627332 453074 627432
rect 453198 627332 453298 627432
rect 453422 627332 453522 627432
rect 453646 627332 453746 627432
rect 453870 627332 453970 627432
rect 454094 627332 454194 627432
rect 454318 627332 454418 627432
rect 454542 627332 454642 627432
rect 454766 627332 454866 627432
rect 454990 627332 455090 627432
rect 455214 627332 455314 627432
rect 455438 627332 455538 627432
rect 455662 627332 455762 627432
rect 455886 627332 455986 627432
rect 449390 627108 449490 627208
rect 449614 627108 449714 627208
rect 449838 627108 449938 627208
rect 450062 627108 450162 627208
rect 450286 627108 450386 627208
rect 450510 627108 450610 627208
rect 450734 627108 450834 627208
rect 450958 627108 451058 627208
rect 451182 627108 451282 627208
rect 451406 627108 451506 627208
rect 451630 627108 451730 627208
rect 451854 627108 451954 627208
rect 452078 627108 452178 627208
rect 452302 627108 452402 627208
rect 452526 627108 452626 627208
rect 452750 627108 452850 627208
rect 452974 627108 453074 627208
rect 453198 627108 453298 627208
rect 453422 627108 453522 627208
rect 453646 627108 453746 627208
rect 453870 627108 453970 627208
rect 454094 627108 454194 627208
rect 454318 627108 454418 627208
rect 454542 627108 454642 627208
rect 454766 627108 454866 627208
rect 454990 627108 455090 627208
rect 455214 627108 455314 627208
rect 455438 627108 455538 627208
rect 455662 627108 455762 627208
rect 455886 627108 455986 627208
rect 449390 626884 449490 626984
rect 449614 626884 449714 626984
rect 449838 626884 449938 626984
rect 450062 626884 450162 626984
rect 450286 626884 450386 626984
rect 450510 626884 450610 626984
rect 450734 626884 450834 626984
rect 450958 626884 451058 626984
rect 451182 626884 451282 626984
rect 451406 626884 451506 626984
rect 451630 626884 451730 626984
rect 451854 626884 451954 626984
rect 452078 626884 452178 626984
rect 452302 626884 452402 626984
rect 452526 626884 452626 626984
rect 452750 626884 452850 626984
rect 452974 626884 453074 626984
rect 453198 626884 453298 626984
rect 453422 626884 453522 626984
rect 453646 626884 453746 626984
rect 453870 626884 453970 626984
rect 454094 626884 454194 626984
rect 454318 626884 454418 626984
rect 454542 626884 454642 626984
rect 454766 626884 454866 626984
rect 454990 626884 455090 626984
rect 455214 626884 455314 626984
rect 455438 626884 455538 626984
rect 455662 626884 455762 626984
rect 455886 626884 455986 626984
rect 449390 626660 449490 626760
rect 449614 626660 449714 626760
rect 449838 626660 449938 626760
rect 450062 626660 450162 626760
rect 450286 626660 450386 626760
rect 450510 626660 450610 626760
rect 450734 626660 450834 626760
rect 450958 626660 451058 626760
rect 451182 626660 451282 626760
rect 451406 626660 451506 626760
rect 451630 626660 451730 626760
rect 451854 626660 451954 626760
rect 452078 626660 452178 626760
rect 452302 626660 452402 626760
rect 452526 626660 452626 626760
rect 452750 626660 452850 626760
rect 452974 626660 453074 626760
rect 453198 626660 453298 626760
rect 453422 626660 453522 626760
rect 453646 626660 453746 626760
rect 453870 626660 453970 626760
rect 454094 626660 454194 626760
rect 454318 626660 454418 626760
rect 454542 626660 454642 626760
rect 454766 626660 454866 626760
rect 454990 626660 455090 626760
rect 455214 626660 455314 626760
rect 455438 626660 455538 626760
rect 455662 626660 455762 626760
rect 455886 626660 455986 626760
rect 475660 627576 475760 627676
rect 475884 627576 475984 627676
rect 476108 627576 476208 627676
rect 476332 627576 476432 627676
rect 476556 627576 476656 627676
rect 476780 627576 476880 627676
rect 477004 627576 477104 627676
rect 477228 627576 477328 627676
rect 477452 627576 477552 627676
rect 477676 627576 477776 627676
rect 477900 627576 478000 627676
rect 478124 627576 478224 627676
rect 478348 627576 478448 627676
rect 478572 627576 478672 627676
rect 478796 627576 478896 627676
rect 479020 627576 479120 627676
rect 479244 627576 479344 627676
rect 479468 627576 479568 627676
rect 479692 627576 479792 627676
rect 479916 627576 480016 627676
rect 480140 627576 480240 627676
rect 480364 627576 480464 627676
rect 480588 627576 480688 627676
rect 480812 627576 480912 627676
rect 481036 627576 481136 627676
rect 481260 627576 481360 627676
rect 481484 627576 481584 627676
rect 481708 627576 481808 627676
rect 481932 627576 482032 627676
rect 482156 627576 482256 627676
rect 475660 627352 475760 627452
rect 475884 627352 475984 627452
rect 476108 627352 476208 627452
rect 476332 627352 476432 627452
rect 476556 627352 476656 627452
rect 476780 627352 476880 627452
rect 477004 627352 477104 627452
rect 477228 627352 477328 627452
rect 477452 627352 477552 627452
rect 477676 627352 477776 627452
rect 477900 627352 478000 627452
rect 478124 627352 478224 627452
rect 478348 627352 478448 627452
rect 478572 627352 478672 627452
rect 478796 627352 478896 627452
rect 479020 627352 479120 627452
rect 479244 627352 479344 627452
rect 479468 627352 479568 627452
rect 479692 627352 479792 627452
rect 479916 627352 480016 627452
rect 480140 627352 480240 627452
rect 480364 627352 480464 627452
rect 480588 627352 480688 627452
rect 480812 627352 480912 627452
rect 481036 627352 481136 627452
rect 481260 627352 481360 627452
rect 481484 627352 481584 627452
rect 481708 627352 481808 627452
rect 481932 627352 482032 627452
rect 482156 627352 482256 627452
rect 475660 627128 475760 627228
rect 475884 627128 475984 627228
rect 476108 627128 476208 627228
rect 476332 627128 476432 627228
rect 476556 627128 476656 627228
rect 476780 627128 476880 627228
rect 477004 627128 477104 627228
rect 477228 627128 477328 627228
rect 477452 627128 477552 627228
rect 477676 627128 477776 627228
rect 477900 627128 478000 627228
rect 478124 627128 478224 627228
rect 478348 627128 478448 627228
rect 478572 627128 478672 627228
rect 478796 627128 478896 627228
rect 479020 627128 479120 627228
rect 479244 627128 479344 627228
rect 479468 627128 479568 627228
rect 479692 627128 479792 627228
rect 479916 627128 480016 627228
rect 480140 627128 480240 627228
rect 480364 627128 480464 627228
rect 480588 627128 480688 627228
rect 480812 627128 480912 627228
rect 481036 627128 481136 627228
rect 481260 627128 481360 627228
rect 481484 627128 481584 627228
rect 481708 627128 481808 627228
rect 481932 627128 482032 627228
rect 482156 627128 482256 627228
rect 475660 626904 475760 627004
rect 475884 626904 475984 627004
rect 476108 626904 476208 627004
rect 476332 626904 476432 627004
rect 476556 626904 476656 627004
rect 476780 626904 476880 627004
rect 477004 626904 477104 627004
rect 477228 626904 477328 627004
rect 477452 626904 477552 627004
rect 477676 626904 477776 627004
rect 477900 626904 478000 627004
rect 478124 626904 478224 627004
rect 478348 626904 478448 627004
rect 478572 626904 478672 627004
rect 478796 626904 478896 627004
rect 479020 626904 479120 627004
rect 479244 626904 479344 627004
rect 479468 626904 479568 627004
rect 479692 626904 479792 627004
rect 479916 626904 480016 627004
rect 480140 626904 480240 627004
rect 480364 626904 480464 627004
rect 480588 626904 480688 627004
rect 480812 626904 480912 627004
rect 481036 626904 481136 627004
rect 481260 626904 481360 627004
rect 481484 626904 481584 627004
rect 481708 626904 481808 627004
rect 481932 626904 482032 627004
rect 482156 626904 482256 627004
rect 475660 626680 475760 626780
rect 475884 626680 475984 626780
rect 476108 626680 476208 626780
rect 476332 626680 476432 626780
rect 476556 626680 476656 626780
rect 476780 626680 476880 626780
rect 477004 626680 477104 626780
rect 477228 626680 477328 626780
rect 477452 626680 477552 626780
rect 477676 626680 477776 626780
rect 477900 626680 478000 626780
rect 478124 626680 478224 626780
rect 478348 626680 478448 626780
rect 478572 626680 478672 626780
rect 478796 626680 478896 626780
rect 479020 626680 479120 626780
rect 479244 626680 479344 626780
rect 479468 626680 479568 626780
rect 479692 626680 479792 626780
rect 479916 626680 480016 626780
rect 480140 626680 480240 626780
rect 480364 626680 480464 626780
rect 480588 626680 480688 626780
rect 480812 626680 480912 626780
rect 481036 626680 481136 626780
rect 481260 626680 481360 626780
rect 481484 626680 481584 626780
rect 481708 626680 481808 626780
rect 481932 626680 482032 626780
rect 482156 626680 482256 626780
<< metal3 >>
rect 428964 662766 435620 669400
rect 459044 668964 474444 669400
rect 428964 657022 429964 662766
rect 434748 657022 435620 662766
rect 428964 649366 435620 657022
rect 438864 662766 456024 663582
rect 438864 657022 438964 662766
rect 443748 657022 444964 662766
rect 449748 657022 450964 662766
rect 455748 657022 456024 662766
rect 459038 662382 474444 668964
rect 438864 654876 456024 657022
rect 438864 654776 438920 654876
rect 439020 654776 439144 654876
rect 439244 654776 439368 654876
rect 439468 654776 439592 654876
rect 439692 654776 439816 654876
rect 439916 654776 440040 654876
rect 440140 654776 440264 654876
rect 440364 654776 440488 654876
rect 440588 654776 440712 654876
rect 440812 654776 440936 654876
rect 441036 654776 441160 654876
rect 441260 654776 441384 654876
rect 441484 654776 441608 654876
rect 441708 654776 441832 654876
rect 441932 654776 442056 654876
rect 442156 654776 442280 654876
rect 442380 654776 442504 654876
rect 442604 654776 442728 654876
rect 442828 654776 442952 654876
rect 443052 654776 443176 654876
rect 443276 654776 443400 654876
rect 443500 654776 443624 654876
rect 443724 654776 443848 654876
rect 443948 654776 444072 654876
rect 444172 654776 444296 654876
rect 444396 654776 444520 654876
rect 444620 654776 444744 654876
rect 444844 654776 444968 654876
rect 445068 654776 445192 654876
rect 445292 654776 445416 654876
rect 445516 654776 449390 654876
rect 449490 654776 449614 654876
rect 449714 654776 449838 654876
rect 449938 654776 450062 654876
rect 450162 654776 450286 654876
rect 450386 654776 450510 654876
rect 450610 654776 450734 654876
rect 450834 654776 450958 654876
rect 451058 654776 451182 654876
rect 451282 654776 451406 654876
rect 451506 654776 451630 654876
rect 451730 654776 451854 654876
rect 451954 654776 452078 654876
rect 452178 654776 452302 654876
rect 452402 654776 452526 654876
rect 452626 654776 452750 654876
rect 452850 654776 452974 654876
rect 453074 654776 453198 654876
rect 453298 654776 453422 654876
rect 453522 654776 453646 654876
rect 453746 654776 453870 654876
rect 453970 654776 454094 654876
rect 454194 654776 454318 654876
rect 454418 654776 454542 654876
rect 454642 654776 454766 654876
rect 454866 654776 454990 654876
rect 455090 654776 455214 654876
rect 455314 654776 455438 654876
rect 455538 654776 455662 654876
rect 455762 654776 455886 654876
rect 455986 654776 456024 654876
rect 438864 654652 456024 654776
rect 438864 654552 438920 654652
rect 439020 654552 439144 654652
rect 439244 654552 439368 654652
rect 439468 654552 439592 654652
rect 439692 654552 439816 654652
rect 439916 654552 440040 654652
rect 440140 654552 440264 654652
rect 440364 654552 440488 654652
rect 440588 654552 440712 654652
rect 440812 654552 440936 654652
rect 441036 654552 441160 654652
rect 441260 654552 441384 654652
rect 441484 654552 441608 654652
rect 441708 654552 441832 654652
rect 441932 654552 442056 654652
rect 442156 654552 442280 654652
rect 442380 654552 442504 654652
rect 442604 654552 442728 654652
rect 442828 654552 442952 654652
rect 443052 654552 443176 654652
rect 443276 654552 443400 654652
rect 443500 654552 443624 654652
rect 443724 654552 443848 654652
rect 443948 654552 444072 654652
rect 444172 654552 444296 654652
rect 444396 654552 444520 654652
rect 444620 654552 444744 654652
rect 444844 654552 444968 654652
rect 445068 654552 445192 654652
rect 445292 654552 445416 654652
rect 445516 654552 449390 654652
rect 449490 654552 449614 654652
rect 449714 654552 449838 654652
rect 449938 654552 450062 654652
rect 450162 654552 450286 654652
rect 450386 654552 450510 654652
rect 450610 654552 450734 654652
rect 450834 654552 450958 654652
rect 451058 654552 451182 654652
rect 451282 654552 451406 654652
rect 451506 654552 451630 654652
rect 451730 654552 451854 654652
rect 451954 654552 452078 654652
rect 452178 654552 452302 654652
rect 452402 654552 452526 654652
rect 452626 654552 452750 654652
rect 452850 654552 452974 654652
rect 453074 654552 453198 654652
rect 453298 654552 453422 654652
rect 453522 654552 453646 654652
rect 453746 654552 453870 654652
rect 453970 654552 454094 654652
rect 454194 654552 454318 654652
rect 454418 654552 454542 654652
rect 454642 654552 454766 654652
rect 454866 654552 454990 654652
rect 455090 654552 455214 654652
rect 455314 654552 455438 654652
rect 455538 654552 455662 654652
rect 455762 654552 455886 654652
rect 455986 654552 456024 654652
rect 438864 654428 456024 654552
rect 438864 654328 438920 654428
rect 439020 654328 439144 654428
rect 439244 654328 439368 654428
rect 439468 654328 439592 654428
rect 439692 654328 439816 654428
rect 439916 654328 440040 654428
rect 440140 654328 440264 654428
rect 440364 654328 440488 654428
rect 440588 654328 440712 654428
rect 440812 654328 440936 654428
rect 441036 654328 441160 654428
rect 441260 654328 441384 654428
rect 441484 654328 441608 654428
rect 441708 654328 441832 654428
rect 441932 654328 442056 654428
rect 442156 654328 442280 654428
rect 442380 654328 442504 654428
rect 442604 654328 442728 654428
rect 442828 654328 442952 654428
rect 443052 654328 443176 654428
rect 443276 654328 443400 654428
rect 443500 654328 443624 654428
rect 443724 654328 443848 654428
rect 443948 654328 444072 654428
rect 444172 654328 444296 654428
rect 444396 654328 444520 654428
rect 444620 654328 444744 654428
rect 444844 654328 444968 654428
rect 445068 654328 445192 654428
rect 445292 654328 445416 654428
rect 445516 654328 449390 654428
rect 449490 654328 449614 654428
rect 449714 654328 449838 654428
rect 449938 654328 450062 654428
rect 450162 654328 450286 654428
rect 450386 654328 450510 654428
rect 450610 654328 450734 654428
rect 450834 654328 450958 654428
rect 451058 654328 451182 654428
rect 451282 654328 451406 654428
rect 451506 654328 451630 654428
rect 451730 654328 451854 654428
rect 451954 654328 452078 654428
rect 452178 654328 452302 654428
rect 452402 654328 452526 654428
rect 452626 654328 452750 654428
rect 452850 654328 452974 654428
rect 453074 654328 453198 654428
rect 453298 654328 453422 654428
rect 453522 654328 453646 654428
rect 453746 654328 453870 654428
rect 453970 654328 454094 654428
rect 454194 654328 454318 654428
rect 454418 654328 454542 654428
rect 454642 654328 454766 654428
rect 454866 654328 454990 654428
rect 455090 654328 455214 654428
rect 455314 654328 455438 654428
rect 455538 654328 455662 654428
rect 455762 654328 455886 654428
rect 455986 654328 456024 654428
rect 438864 654204 456024 654328
rect 438864 654104 438920 654204
rect 439020 654104 439144 654204
rect 439244 654104 439368 654204
rect 439468 654104 439592 654204
rect 439692 654104 439816 654204
rect 439916 654104 440040 654204
rect 440140 654104 440264 654204
rect 440364 654104 440488 654204
rect 440588 654104 440712 654204
rect 440812 654104 440936 654204
rect 441036 654104 441160 654204
rect 441260 654104 441384 654204
rect 441484 654104 441608 654204
rect 441708 654104 441832 654204
rect 441932 654104 442056 654204
rect 442156 654104 442280 654204
rect 442380 654104 442504 654204
rect 442604 654104 442728 654204
rect 442828 654104 442952 654204
rect 443052 654104 443176 654204
rect 443276 654104 443400 654204
rect 443500 654104 443624 654204
rect 443724 654104 443848 654204
rect 443948 654104 444072 654204
rect 444172 654104 444296 654204
rect 444396 654104 444520 654204
rect 444620 654104 444744 654204
rect 444844 654104 444968 654204
rect 445068 654104 445192 654204
rect 445292 654104 445416 654204
rect 445516 654104 449390 654204
rect 449490 654104 449614 654204
rect 449714 654104 449838 654204
rect 449938 654104 450062 654204
rect 450162 654104 450286 654204
rect 450386 654104 450510 654204
rect 450610 654104 450734 654204
rect 450834 654104 450958 654204
rect 451058 654104 451182 654204
rect 451282 654104 451406 654204
rect 451506 654104 451630 654204
rect 451730 654104 451854 654204
rect 451954 654104 452078 654204
rect 452178 654104 452302 654204
rect 452402 654104 452526 654204
rect 452626 654104 452750 654204
rect 452850 654104 452974 654204
rect 453074 654104 453198 654204
rect 453298 654104 453422 654204
rect 453522 654104 453646 654204
rect 453746 654104 453870 654204
rect 453970 654104 454094 654204
rect 454194 654104 454318 654204
rect 454418 654104 454542 654204
rect 454642 654104 454766 654204
rect 454866 654104 454990 654204
rect 455090 654104 455214 654204
rect 455314 654104 455438 654204
rect 455538 654104 455662 654204
rect 455762 654104 455886 654204
rect 455986 654104 456024 654204
rect 438864 653980 456024 654104
rect 438864 653880 438920 653980
rect 439020 653880 439144 653980
rect 439244 653880 439368 653980
rect 439468 653880 439592 653980
rect 439692 653880 439816 653980
rect 439916 653880 440040 653980
rect 440140 653880 440264 653980
rect 440364 653880 440488 653980
rect 440588 653880 440712 653980
rect 440812 653880 440936 653980
rect 441036 653880 441160 653980
rect 441260 653880 441384 653980
rect 441484 653880 441608 653980
rect 441708 653880 441832 653980
rect 441932 653880 442056 653980
rect 442156 653880 442280 653980
rect 442380 653880 442504 653980
rect 442604 653880 442728 653980
rect 442828 653880 442952 653980
rect 443052 653880 443176 653980
rect 443276 653880 443400 653980
rect 443500 653880 443624 653980
rect 443724 653880 443848 653980
rect 443948 653880 444072 653980
rect 444172 653880 444296 653980
rect 444396 653880 444520 653980
rect 444620 653880 444744 653980
rect 444844 653880 444968 653980
rect 445068 653880 445192 653980
rect 445292 653880 445416 653980
rect 445516 653880 449390 653980
rect 449490 653880 449614 653980
rect 449714 653880 449838 653980
rect 449938 653880 450062 653980
rect 450162 653880 450286 653980
rect 450386 653880 450510 653980
rect 450610 653880 450734 653980
rect 450834 653880 450958 653980
rect 451058 653880 451182 653980
rect 451282 653880 451406 653980
rect 451506 653880 451630 653980
rect 451730 653880 451854 653980
rect 451954 653880 452078 653980
rect 452178 653880 452302 653980
rect 452402 653880 452526 653980
rect 452626 653880 452750 653980
rect 452850 653880 452974 653980
rect 453074 653880 453198 653980
rect 453298 653880 453422 653980
rect 453522 653880 453646 653980
rect 453746 653880 453870 653980
rect 453970 653880 454094 653980
rect 454194 653880 454318 653980
rect 454418 653880 454542 653980
rect 454642 653880 454766 653980
rect 454866 653880 454990 653980
rect 455090 653880 455214 653980
rect 455314 653880 455438 653980
rect 455538 653880 455662 653980
rect 455762 653880 455886 653980
rect 455986 653880 456024 653980
rect 438864 653842 456024 653880
rect 440681 652769 451967 652775
rect 440681 651913 440687 652769
rect 451961 651913 451967 652769
rect 440681 651907 451967 651913
rect 428964 643622 429964 649366
rect 434748 643622 435620 649366
rect 428964 635966 435620 643622
rect 437864 650178 438924 650202
rect 437864 650078 437894 650178
rect 437994 650078 438118 650178
rect 438218 650078 438342 650178
rect 438442 650078 438566 650178
rect 438666 650078 438790 650178
rect 438890 650078 438924 650178
rect 437864 649954 438924 650078
rect 437864 649854 437894 649954
rect 437994 649854 438118 649954
rect 438218 649854 438342 649954
rect 438442 649854 438566 649954
rect 438666 649854 438790 649954
rect 438890 649854 438924 649954
rect 437864 649730 438924 649854
rect 437864 649630 437894 649730
rect 437994 649630 438118 649730
rect 438218 649630 438342 649730
rect 438442 649630 438566 649730
rect 438666 649630 438790 649730
rect 438890 649630 438924 649730
rect 437864 649506 438924 649630
rect 437864 649406 437894 649506
rect 437994 649406 438118 649506
rect 438218 649406 438342 649506
rect 438442 649406 438566 649506
rect 438666 649406 438790 649506
rect 438890 649406 438924 649506
rect 437864 649282 438924 649406
rect 437864 649182 437894 649282
rect 437994 649182 438118 649282
rect 438218 649182 438342 649282
rect 438442 649182 438566 649282
rect 438666 649182 438790 649282
rect 438890 649182 438924 649282
rect 437864 649058 438924 649182
rect 437864 648958 437894 649058
rect 437994 648958 438118 649058
rect 438218 648958 438342 649058
rect 438442 648958 438566 649058
rect 438666 648958 438790 649058
rect 438890 648958 438924 649058
rect 437864 648834 438924 648958
rect 437864 648734 437894 648834
rect 437994 648734 438118 648834
rect 438218 648734 438342 648834
rect 438442 648734 438566 648834
rect 438666 648734 438790 648834
rect 438890 648734 438924 648834
rect 437864 648610 438924 648734
rect 437864 648510 437894 648610
rect 437994 648510 438118 648610
rect 438218 648510 438342 648610
rect 438442 648510 438566 648610
rect 438666 648510 438790 648610
rect 438890 648510 438924 648610
rect 437864 648386 438924 648510
rect 437864 648286 437894 648386
rect 437994 648286 438118 648386
rect 438218 648286 438342 648386
rect 438442 648286 438566 648386
rect 438666 648286 438790 648386
rect 438890 648286 438924 648386
rect 437864 648162 438924 648286
rect 437864 648062 437894 648162
rect 437994 648062 438118 648162
rect 438218 648062 438342 648162
rect 438442 648062 438566 648162
rect 438666 648062 438790 648162
rect 438890 648062 438924 648162
rect 437864 647938 438924 648062
rect 437864 647838 437894 647938
rect 437994 647838 438118 647938
rect 438218 647838 438342 647938
rect 438442 647838 438566 647938
rect 438666 647838 438790 647938
rect 438890 647838 438924 647938
rect 437864 647714 438924 647838
rect 437864 647614 437894 647714
rect 437994 647614 438118 647714
rect 438218 647614 438342 647714
rect 438442 647614 438566 647714
rect 438666 647614 438790 647714
rect 438890 647614 438924 647714
rect 437864 647490 438924 647614
rect 437864 647390 437894 647490
rect 437994 647390 438118 647490
rect 438218 647390 438342 647490
rect 438442 647390 438566 647490
rect 438666 647390 438790 647490
rect 438890 647390 438924 647490
rect 437864 647266 438924 647390
rect 437864 647166 437894 647266
rect 437994 647166 438118 647266
rect 438218 647166 438342 647266
rect 438442 647166 438566 647266
rect 438666 647166 438790 647266
rect 438890 647166 438924 647266
rect 437864 647042 438924 647166
rect 437864 646942 437894 647042
rect 437994 646942 438118 647042
rect 438218 646942 438342 647042
rect 438442 646942 438566 647042
rect 438666 646942 438790 647042
rect 438890 646942 438924 647042
rect 437864 646818 438924 646942
rect 437864 646718 437894 646818
rect 437994 646718 438118 646818
rect 438218 646718 438342 646818
rect 438442 646718 438566 646818
rect 438666 646718 438790 646818
rect 438890 646718 438924 646818
rect 437864 646594 438924 646718
rect 437864 646494 437894 646594
rect 437994 646494 438118 646594
rect 438218 646494 438342 646594
rect 438442 646494 438566 646594
rect 438666 646494 438790 646594
rect 438890 646494 438924 646594
rect 437864 646370 438924 646494
rect 437864 646270 437894 646370
rect 437994 646270 438118 646370
rect 438218 646270 438342 646370
rect 438442 646270 438566 646370
rect 438666 646270 438790 646370
rect 438890 646270 438924 646370
rect 437864 646146 438924 646270
rect 437864 646046 437894 646146
rect 437994 646046 438118 646146
rect 438218 646046 438342 646146
rect 438442 646046 438566 646146
rect 438666 646046 438790 646146
rect 438890 646046 438924 646146
rect 437864 645922 438924 646046
rect 437864 645822 437894 645922
rect 437994 645822 438118 645922
rect 438218 645822 438342 645922
rect 438442 645822 438566 645922
rect 438666 645822 438790 645922
rect 438890 645822 438924 645922
rect 437864 645698 438924 645822
rect 437864 645598 437894 645698
rect 437994 645598 438118 645698
rect 438218 645598 438342 645698
rect 438442 645598 438566 645698
rect 438666 645598 438790 645698
rect 438890 645598 438924 645698
rect 437864 645474 438924 645598
rect 437864 645374 437894 645474
rect 437994 645374 438118 645474
rect 438218 645374 438342 645474
rect 438442 645374 438566 645474
rect 438666 645374 438790 645474
rect 438890 645374 438924 645474
rect 437864 645250 438924 645374
rect 437864 645150 437894 645250
rect 437994 645150 438118 645250
rect 438218 645150 438342 645250
rect 438442 645150 438566 645250
rect 438666 645150 438790 645250
rect 438890 645150 438924 645250
rect 437864 645026 438924 645150
rect 437864 644926 437894 645026
rect 437994 644926 438118 645026
rect 438218 644926 438342 645026
rect 438442 644926 438566 645026
rect 438666 644926 438790 645026
rect 438890 644926 438924 645026
rect 437864 644802 438924 644926
rect 437864 644702 437894 644802
rect 437994 644702 438118 644802
rect 438218 644702 438342 644802
rect 438442 644702 438566 644802
rect 438666 644702 438790 644802
rect 438890 644702 438924 644802
rect 437864 644578 438924 644702
rect 437864 644478 437894 644578
rect 437994 644478 438118 644578
rect 438218 644478 438342 644578
rect 438442 644478 438566 644578
rect 438666 644478 438790 644578
rect 438890 644478 438924 644578
rect 437864 644354 438924 644478
rect 437864 644254 437894 644354
rect 437994 644254 438118 644354
rect 438218 644254 438342 644354
rect 438442 644254 438566 644354
rect 438666 644254 438790 644354
rect 438890 644254 438924 644354
rect 437864 644130 438924 644254
rect 437864 644030 437894 644130
rect 437994 644030 438118 644130
rect 438218 644030 438342 644130
rect 438442 644030 438566 644130
rect 438666 644030 438790 644130
rect 438890 644030 438924 644130
rect 437864 643906 438924 644030
rect 437864 643806 437894 643906
rect 437994 643806 438118 643906
rect 438218 643806 438342 643906
rect 438442 643806 438566 643906
rect 438666 643806 438790 643906
rect 438890 643806 438924 643906
rect 437864 643682 438924 643806
rect 437864 643582 437894 643682
rect 437994 643582 438118 643682
rect 438218 643582 438342 643682
rect 438442 643582 438566 643682
rect 438666 643582 438790 643682
rect 438890 643582 438924 643682
rect 437864 643542 438924 643582
rect 444360 644326 451530 644354
rect 444360 643782 444975 644326
rect 445039 643782 445694 644326
rect 445758 643782 446413 644326
rect 446477 643782 447132 644326
rect 447196 643782 447851 644326
rect 447915 643782 448570 644326
rect 448634 643782 449289 644326
rect 449353 643782 450008 644326
rect 450072 643782 450727 644326
rect 450791 643782 451446 644326
rect 451510 643782 451530 644326
rect 444360 643626 451530 643782
rect 444360 643082 444975 643626
rect 445039 643082 445694 643626
rect 445758 643082 446413 643626
rect 446477 643082 447132 643626
rect 447196 643082 447851 643626
rect 447915 643082 448570 643626
rect 448634 643082 449289 643626
rect 449353 643082 450008 643626
rect 450072 643082 450727 643626
rect 450791 643082 451446 643626
rect 451510 643082 451530 643626
rect 444360 642926 451530 643082
rect 444360 642382 444975 642926
rect 445039 642382 445694 642926
rect 445758 642382 446413 642926
rect 446477 642382 447132 642926
rect 447196 642382 447851 642926
rect 447915 642382 448570 642926
rect 448634 642382 449289 642926
rect 449353 642382 450008 642926
rect 450072 642382 450727 642926
rect 450791 642382 451446 642926
rect 451510 642382 451530 642926
rect 444360 642226 451530 642382
rect 444360 641682 444975 642226
rect 445039 641682 445694 642226
rect 445758 641682 446413 642226
rect 446477 641682 447132 642226
rect 447196 641682 447851 642226
rect 447915 641682 448570 642226
rect 448634 641682 449289 642226
rect 449353 641682 450008 642226
rect 450072 641682 450727 642226
rect 450791 641682 451446 642226
rect 451510 641682 451530 642226
rect 444360 641526 451530 641682
rect 444360 640982 444975 641526
rect 445039 640982 445694 641526
rect 445758 640982 446413 641526
rect 446477 640982 447132 641526
rect 447196 640982 447851 641526
rect 447915 640982 448570 641526
rect 448634 640982 449289 641526
rect 449353 640982 450008 641526
rect 450072 640982 450727 641526
rect 450791 640982 451446 641526
rect 451510 640982 451530 641526
rect 444360 640826 451530 640982
rect 444360 640282 444975 640826
rect 445039 640282 445694 640826
rect 445758 640282 446413 640826
rect 446477 640282 447132 640826
rect 447196 640282 447851 640826
rect 447915 640282 448570 640826
rect 448634 640282 449289 640826
rect 449353 640282 450008 640826
rect 450072 640282 450727 640826
rect 450791 640282 451446 640826
rect 451510 640282 451530 640826
rect 444360 640126 451530 640282
rect 444360 639582 444975 640126
rect 445039 639582 445694 640126
rect 445758 639582 446413 640126
rect 446477 639582 447132 640126
rect 447196 639582 447851 640126
rect 447915 639582 448570 640126
rect 448634 639582 449289 640126
rect 449353 639582 450008 640126
rect 450072 639582 450727 640126
rect 450791 639582 451446 640126
rect 451510 639582 451530 640126
rect 459044 641050 474444 662382
rect 475624 663086 482444 663562
rect 475624 657342 476524 663086
rect 481308 657342 482444 663086
rect 475624 654926 482444 657342
rect 475620 654896 482444 654926
rect 475620 654796 475660 654896
rect 475760 654796 475884 654896
rect 475984 654796 476108 654896
rect 476208 654796 476332 654896
rect 476432 654796 476556 654896
rect 476656 654796 476780 654896
rect 476880 654796 477004 654896
rect 477104 654796 477228 654896
rect 477328 654796 477452 654896
rect 477552 654796 477676 654896
rect 477776 654796 477900 654896
rect 478000 654796 478124 654896
rect 478224 654796 478348 654896
rect 478448 654796 478572 654896
rect 478672 654796 478796 654896
rect 478896 654796 479020 654896
rect 479120 654796 479244 654896
rect 479344 654796 479468 654896
rect 479568 654796 479692 654896
rect 479792 654796 479916 654896
rect 480016 654796 480140 654896
rect 480240 654796 480364 654896
rect 480464 654796 480588 654896
rect 480688 654796 480812 654896
rect 480912 654796 481036 654896
rect 481136 654796 481260 654896
rect 481360 654796 481484 654896
rect 481584 654796 481708 654896
rect 481808 654796 481932 654896
rect 482032 654796 482156 654896
rect 482256 654796 482444 654896
rect 475620 654672 482444 654796
rect 475620 654572 475660 654672
rect 475760 654572 475884 654672
rect 475984 654572 476108 654672
rect 476208 654572 476332 654672
rect 476432 654572 476556 654672
rect 476656 654572 476780 654672
rect 476880 654572 477004 654672
rect 477104 654572 477228 654672
rect 477328 654572 477452 654672
rect 477552 654572 477676 654672
rect 477776 654572 477900 654672
rect 478000 654572 478124 654672
rect 478224 654572 478348 654672
rect 478448 654572 478572 654672
rect 478672 654572 478796 654672
rect 478896 654572 479020 654672
rect 479120 654572 479244 654672
rect 479344 654572 479468 654672
rect 479568 654572 479692 654672
rect 479792 654572 479916 654672
rect 480016 654572 480140 654672
rect 480240 654572 480364 654672
rect 480464 654572 480588 654672
rect 480688 654572 480812 654672
rect 480912 654572 481036 654672
rect 481136 654572 481260 654672
rect 481360 654572 481484 654672
rect 481584 654572 481708 654672
rect 481808 654572 481932 654672
rect 482032 654572 482156 654672
rect 482256 654572 482444 654672
rect 475620 654448 482444 654572
rect 475620 654348 475660 654448
rect 475760 654348 475884 654448
rect 475984 654348 476108 654448
rect 476208 654348 476332 654448
rect 476432 654348 476556 654448
rect 476656 654348 476780 654448
rect 476880 654348 477004 654448
rect 477104 654348 477228 654448
rect 477328 654348 477452 654448
rect 477552 654348 477676 654448
rect 477776 654348 477900 654448
rect 478000 654348 478124 654448
rect 478224 654348 478348 654448
rect 478448 654348 478572 654448
rect 478672 654348 478796 654448
rect 478896 654348 479020 654448
rect 479120 654348 479244 654448
rect 479344 654348 479468 654448
rect 479568 654348 479692 654448
rect 479792 654348 479916 654448
rect 480016 654348 480140 654448
rect 480240 654348 480364 654448
rect 480464 654348 480588 654448
rect 480688 654348 480812 654448
rect 480912 654348 481036 654448
rect 481136 654348 481260 654448
rect 481360 654348 481484 654448
rect 481584 654348 481708 654448
rect 481808 654348 481932 654448
rect 482032 654348 482156 654448
rect 482256 654348 482444 654448
rect 475620 654224 482444 654348
rect 475620 654124 475660 654224
rect 475760 654124 475884 654224
rect 475984 654124 476108 654224
rect 476208 654124 476332 654224
rect 476432 654124 476556 654224
rect 476656 654124 476780 654224
rect 476880 654124 477004 654224
rect 477104 654124 477228 654224
rect 477328 654124 477452 654224
rect 477552 654124 477676 654224
rect 477776 654124 477900 654224
rect 478000 654124 478124 654224
rect 478224 654124 478348 654224
rect 478448 654124 478572 654224
rect 478672 654124 478796 654224
rect 478896 654124 479020 654224
rect 479120 654124 479244 654224
rect 479344 654124 479468 654224
rect 479568 654124 479692 654224
rect 479792 654124 479916 654224
rect 480016 654124 480140 654224
rect 480240 654124 480364 654224
rect 480464 654124 480588 654224
rect 480688 654124 480812 654224
rect 480912 654124 481036 654224
rect 481136 654124 481260 654224
rect 481360 654124 481484 654224
rect 481584 654124 481708 654224
rect 481808 654124 481932 654224
rect 482032 654124 482156 654224
rect 482256 654124 482444 654224
rect 475620 654000 482444 654124
rect 475620 653900 475660 654000
rect 475760 653900 475884 654000
rect 475984 653900 476108 654000
rect 476208 653900 476332 654000
rect 476432 653900 476556 654000
rect 476656 653900 476780 654000
rect 476880 653900 477004 654000
rect 477104 653900 477228 654000
rect 477328 653900 477452 654000
rect 477552 653900 477676 654000
rect 477776 653900 477900 654000
rect 478000 653900 478124 654000
rect 478224 653900 478348 654000
rect 478448 653900 478572 654000
rect 478672 653900 478796 654000
rect 478896 653900 479020 654000
rect 479120 653900 479244 654000
rect 479344 653900 479468 654000
rect 479568 653900 479692 654000
rect 479792 653900 479916 654000
rect 480016 653900 480140 654000
rect 480240 653900 480364 654000
rect 480464 653900 480588 654000
rect 480688 653900 480812 654000
rect 480912 653900 481036 654000
rect 481136 653900 481260 654000
rect 481360 653900 481484 654000
rect 481584 653900 481708 654000
rect 481808 653900 481932 654000
rect 482032 653900 482156 654000
rect 482256 653900 482444 654000
rect 475620 653866 482444 653900
rect 475624 653842 482444 653866
rect 486272 663144 492928 669400
rect 486272 657400 487200 663144
rect 491984 657400 492928 663144
rect 482144 650178 483204 650202
rect 482144 650078 482174 650178
rect 482274 650078 482398 650178
rect 482498 650078 482622 650178
rect 482722 650078 482846 650178
rect 482946 650078 483070 650178
rect 483170 650078 483204 650178
rect 482144 649954 483204 650078
rect 482144 649854 482174 649954
rect 482274 649854 482398 649954
rect 482498 649854 482622 649954
rect 482722 649854 482846 649954
rect 482946 649854 483070 649954
rect 483170 649854 483204 649954
rect 482144 649730 483204 649854
rect 482144 649630 482174 649730
rect 482274 649630 482398 649730
rect 482498 649630 482622 649730
rect 482722 649630 482846 649730
rect 482946 649630 483070 649730
rect 483170 649630 483204 649730
rect 482144 649506 483204 649630
rect 482144 649406 482174 649506
rect 482274 649406 482398 649506
rect 482498 649406 482622 649506
rect 482722 649406 482846 649506
rect 482946 649406 483070 649506
rect 483170 649406 483204 649506
rect 482144 649282 483204 649406
rect 482144 649182 482174 649282
rect 482274 649182 482398 649282
rect 482498 649182 482622 649282
rect 482722 649182 482846 649282
rect 482946 649182 483070 649282
rect 483170 649182 483204 649282
rect 482144 649058 483204 649182
rect 482144 648958 482174 649058
rect 482274 648958 482398 649058
rect 482498 648958 482622 649058
rect 482722 648958 482846 649058
rect 482946 648958 483070 649058
rect 483170 648958 483204 649058
rect 482144 648834 483204 648958
rect 482144 648734 482174 648834
rect 482274 648734 482398 648834
rect 482498 648734 482622 648834
rect 482722 648734 482846 648834
rect 482946 648734 483070 648834
rect 483170 648734 483204 648834
rect 482144 648610 483204 648734
rect 482144 648510 482174 648610
rect 482274 648510 482398 648610
rect 482498 648510 482622 648610
rect 482722 648510 482846 648610
rect 482946 648510 483070 648610
rect 483170 648510 483204 648610
rect 482144 648386 483204 648510
rect 482144 648286 482174 648386
rect 482274 648286 482398 648386
rect 482498 648286 482622 648386
rect 482722 648286 482846 648386
rect 482946 648286 483070 648386
rect 483170 648286 483204 648386
rect 482144 648162 483204 648286
rect 482144 648062 482174 648162
rect 482274 648062 482398 648162
rect 482498 648062 482622 648162
rect 482722 648062 482846 648162
rect 482946 648062 483070 648162
rect 483170 648062 483204 648162
rect 482144 647938 483204 648062
rect 482144 647838 482174 647938
rect 482274 647838 482398 647938
rect 482498 647838 482622 647938
rect 482722 647838 482846 647938
rect 482946 647838 483070 647938
rect 483170 647838 483204 647938
rect 482144 647714 483204 647838
rect 482144 647614 482174 647714
rect 482274 647614 482398 647714
rect 482498 647614 482622 647714
rect 482722 647614 482846 647714
rect 482946 647614 483070 647714
rect 483170 647614 483204 647714
rect 482144 647490 483204 647614
rect 482144 647390 482174 647490
rect 482274 647390 482398 647490
rect 482498 647390 482622 647490
rect 482722 647390 482846 647490
rect 482946 647390 483070 647490
rect 483170 647390 483204 647490
rect 482144 647266 483204 647390
rect 482144 647166 482174 647266
rect 482274 647166 482398 647266
rect 482498 647166 482622 647266
rect 482722 647166 482846 647266
rect 482946 647166 483070 647266
rect 483170 647166 483204 647266
rect 482144 647042 483204 647166
rect 482144 646942 482174 647042
rect 482274 646942 482398 647042
rect 482498 646942 482622 647042
rect 482722 646942 482846 647042
rect 482946 646942 483070 647042
rect 483170 646942 483204 647042
rect 482144 646818 483204 646942
rect 482144 646718 482174 646818
rect 482274 646718 482398 646818
rect 482498 646718 482622 646818
rect 482722 646718 482846 646818
rect 482946 646718 483070 646818
rect 483170 646718 483204 646818
rect 482144 646594 483204 646718
rect 482144 646494 482174 646594
rect 482274 646494 482398 646594
rect 482498 646494 482622 646594
rect 482722 646494 482846 646594
rect 482946 646494 483070 646594
rect 483170 646494 483204 646594
rect 482144 646370 483204 646494
rect 482144 646270 482174 646370
rect 482274 646270 482398 646370
rect 482498 646270 482622 646370
rect 482722 646270 482846 646370
rect 482946 646270 483070 646370
rect 483170 646270 483204 646370
rect 482144 646146 483204 646270
rect 482144 646046 482174 646146
rect 482274 646046 482398 646146
rect 482498 646046 482622 646146
rect 482722 646046 482846 646146
rect 482946 646046 483070 646146
rect 483170 646046 483204 646146
rect 482144 645922 483204 646046
rect 482144 645822 482174 645922
rect 482274 645822 482398 645922
rect 482498 645822 482622 645922
rect 482722 645822 482846 645922
rect 482946 645822 483070 645922
rect 483170 645822 483204 645922
rect 482144 645698 483204 645822
rect 482144 645598 482174 645698
rect 482274 645598 482398 645698
rect 482498 645598 482622 645698
rect 482722 645598 482846 645698
rect 482946 645598 483070 645698
rect 483170 645598 483204 645698
rect 482144 645474 483204 645598
rect 482144 645374 482174 645474
rect 482274 645374 482398 645474
rect 482498 645374 482622 645474
rect 482722 645374 482846 645474
rect 482946 645374 483070 645474
rect 483170 645374 483204 645474
rect 482144 645250 483204 645374
rect 482144 645150 482174 645250
rect 482274 645150 482398 645250
rect 482498 645150 482622 645250
rect 482722 645150 482846 645250
rect 482946 645150 483070 645250
rect 483170 645150 483204 645250
rect 482144 645026 483204 645150
rect 482144 644926 482174 645026
rect 482274 644926 482398 645026
rect 482498 644926 482622 645026
rect 482722 644926 482846 645026
rect 482946 644926 483070 645026
rect 483170 644926 483204 645026
rect 482144 644802 483204 644926
rect 482144 644702 482174 644802
rect 482274 644702 482398 644802
rect 482498 644702 482622 644802
rect 482722 644702 482846 644802
rect 482946 644702 483070 644802
rect 483170 644702 483204 644802
rect 482144 644578 483204 644702
rect 482144 644478 482174 644578
rect 482274 644478 482398 644578
rect 482498 644478 482622 644578
rect 482722 644478 482846 644578
rect 482946 644478 483070 644578
rect 483170 644478 483204 644578
rect 482144 644354 483204 644478
rect 482144 644254 482174 644354
rect 482274 644254 482398 644354
rect 482498 644254 482622 644354
rect 482722 644254 482846 644354
rect 482946 644254 483070 644354
rect 483170 644254 483204 644354
rect 482144 644130 483204 644254
rect 482144 644030 482174 644130
rect 482274 644030 482398 644130
rect 482498 644030 482622 644130
rect 482722 644030 482846 644130
rect 482946 644030 483070 644130
rect 483170 644030 483204 644130
rect 482144 643906 483204 644030
rect 482144 643806 482174 643906
rect 482274 643806 482398 643906
rect 482498 643806 482622 643906
rect 482722 643806 482846 643906
rect 482946 643806 483070 643906
rect 483170 643806 483204 643906
rect 482144 643682 483204 643806
rect 482144 643582 482174 643682
rect 482274 643582 482398 643682
rect 482498 643582 482622 643682
rect 482722 643582 482846 643682
rect 482946 643582 483070 643682
rect 483170 643582 483204 643682
rect 482144 643542 483204 643582
rect 486272 649744 492928 657400
rect 486272 644000 487200 649744
rect 491984 644000 492928 649744
rect 459044 640850 459444 641050
rect 459644 640850 459878 641050
rect 460078 640850 460312 641050
rect 460512 640850 460746 641050
rect 460946 640850 461180 641050
rect 461380 640850 461614 641050
rect 461814 640850 462048 641050
rect 462248 640850 462482 641050
rect 462682 640850 462916 641050
rect 463116 640850 463350 641050
rect 463550 640850 463784 641050
rect 463984 640850 464184 641050
rect 464384 640850 464584 641050
rect 464784 640850 464984 641050
rect 465184 640850 465384 641050
rect 465584 640850 465784 641050
rect 465984 640850 466184 641050
rect 466384 640850 466584 641050
rect 466784 640850 466984 641050
rect 467184 640850 467384 641050
rect 467584 640850 468984 641050
rect 469184 640850 469384 641050
rect 469584 640850 469784 641050
rect 469984 640850 470184 641050
rect 470384 640850 470584 641050
rect 470784 640850 470984 641050
rect 471184 640850 471384 641050
rect 471584 640850 471784 641050
rect 471984 640850 472184 641050
rect 472384 640850 474444 641050
rect 459044 640616 474444 640850
rect 459044 640416 459444 640616
rect 459644 640416 459878 640616
rect 460078 640416 460312 640616
rect 460512 640416 460746 640616
rect 460946 640416 461180 640616
rect 461380 640416 461614 640616
rect 461814 640416 462048 640616
rect 462248 640416 462482 640616
rect 462682 640416 462916 640616
rect 463116 640416 463350 640616
rect 463550 640416 463784 640616
rect 463984 640416 474444 640616
rect 459044 640182 474444 640416
rect 459044 639982 459444 640182
rect 459644 639982 459878 640182
rect 460078 639982 460312 640182
rect 460512 639982 460746 640182
rect 460946 639982 461180 640182
rect 461380 639982 461614 640182
rect 461814 639982 462048 640182
rect 462248 639982 462482 640182
rect 462682 639982 462916 640182
rect 463116 639982 463350 640182
rect 463550 639982 463784 640182
rect 463984 639982 474444 640182
rect 459044 639782 474444 639982
rect 444360 639426 451530 639582
rect 444360 638882 444975 639426
rect 445039 638882 445694 639426
rect 445758 638882 446413 639426
rect 446477 638882 447132 639426
rect 447196 638882 447851 639426
rect 447915 638882 448570 639426
rect 448634 638882 449289 639426
rect 449353 638882 450008 639426
rect 450072 638882 450727 639426
rect 450791 638882 451446 639426
rect 451510 638882 451530 639426
rect 444360 638726 451530 638882
rect 437836 638358 443596 638422
rect 437836 638294 437900 638358
rect 437964 638294 438028 638358
rect 438092 638294 438156 638358
rect 438220 638294 438284 638358
rect 438348 638294 438412 638358
rect 438476 638294 438540 638358
rect 438604 638294 438668 638358
rect 438732 638294 438796 638358
rect 438860 638294 438924 638358
rect 438988 638294 443596 638358
rect 437836 638230 443596 638294
rect 437836 638166 437900 638230
rect 437964 638166 438028 638230
rect 438092 638166 438156 638230
rect 438220 638166 438284 638230
rect 438348 638166 438412 638230
rect 438476 638166 438540 638230
rect 438604 638166 438668 638230
rect 438732 638166 438796 638230
rect 438860 638166 438924 638230
rect 438988 638212 443596 638230
rect 438988 638166 443024 638212
rect 437836 638152 443024 638166
rect 443084 638152 443144 638212
rect 443204 638152 443264 638212
rect 443324 638152 443384 638212
rect 443444 638152 443504 638212
rect 443564 638152 443596 638212
rect 437836 638102 443596 638152
rect 437836 638038 437900 638102
rect 437964 638038 438028 638102
rect 438092 638038 438156 638102
rect 438220 638038 438284 638102
rect 438348 638038 438412 638102
rect 438476 638038 438540 638102
rect 438604 638038 438668 638102
rect 438732 638038 438796 638102
rect 438860 638038 438924 638102
rect 438988 638092 443596 638102
rect 438988 638038 443024 638092
rect 437836 638032 443024 638038
rect 443084 638032 443144 638092
rect 443204 638032 443264 638092
rect 443324 638032 443384 638092
rect 443444 638032 443504 638092
rect 443564 638032 443596 638092
rect 437836 637974 443596 638032
rect 437836 637910 437900 637974
rect 437964 637910 438028 637974
rect 438092 637910 438156 637974
rect 438220 637910 438284 637974
rect 438348 637910 438412 637974
rect 438476 637910 438540 637974
rect 438604 637910 438668 637974
rect 438732 637910 438796 637974
rect 438860 637910 438924 637974
rect 438988 637910 443596 637974
rect 437836 637846 443596 637910
rect 444360 638182 444975 638726
rect 445039 638182 445694 638726
rect 445758 638182 446413 638726
rect 446477 638182 447132 638726
rect 447196 638182 447851 638726
rect 447915 638182 448570 638726
rect 448634 638182 449289 638726
rect 449353 638182 450008 638726
rect 450072 638182 450727 638726
rect 450791 638182 451446 638726
rect 451510 638182 451530 638726
rect 452991 639474 473323 639479
rect 452991 638490 452996 639474
rect 473318 638490 473323 639474
rect 452991 638485 473323 638490
rect 444360 638026 451530 638182
rect 444360 637482 444975 638026
rect 445039 637482 445694 638026
rect 445758 637482 446413 638026
rect 446477 637482 447132 638026
rect 447196 637482 447851 638026
rect 447915 637482 448570 638026
rect 448634 637482 449289 638026
rect 449353 637482 450008 638026
rect 450072 637482 450727 638026
rect 450791 637482 451446 638026
rect 451510 637482 451530 638026
rect 437864 636782 438922 636788
rect 428964 630222 429964 635966
rect 434748 630222 435620 635966
rect 428964 622946 435620 630222
rect 437764 636778 438924 636782
rect 437764 636678 437894 636778
rect 437994 636678 438118 636778
rect 438218 636678 438342 636778
rect 438442 636678 438566 636778
rect 438666 636678 438790 636778
rect 438890 636678 438924 636778
rect 437764 636554 438924 636678
rect 437764 636454 437894 636554
rect 437994 636454 438118 636554
rect 438218 636454 438342 636554
rect 438442 636454 438566 636554
rect 438666 636454 438790 636554
rect 438890 636454 438924 636554
rect 437764 636330 438924 636454
rect 437764 636230 437894 636330
rect 437994 636230 438118 636330
rect 438218 636230 438342 636330
rect 438442 636230 438566 636330
rect 438666 636230 438790 636330
rect 438890 636230 438924 636330
rect 437764 636106 438924 636230
rect 437764 636006 437894 636106
rect 437994 636006 438118 636106
rect 438218 636006 438342 636106
rect 438442 636006 438566 636106
rect 438666 636006 438790 636106
rect 438890 636006 438924 636106
rect 437764 635882 438924 636006
rect 437764 635782 437894 635882
rect 437994 635782 438118 635882
rect 438218 635782 438342 635882
rect 438442 635782 438566 635882
rect 438666 635782 438790 635882
rect 438890 635782 438924 635882
rect 437764 635658 438924 635782
rect 437764 635558 437894 635658
rect 437994 635558 438118 635658
rect 438218 635558 438342 635658
rect 438442 635558 438566 635658
rect 438666 635558 438790 635658
rect 438890 635558 438924 635658
rect 437764 635434 438924 635558
rect 437764 635334 437894 635434
rect 437994 635334 438118 635434
rect 438218 635334 438342 635434
rect 438442 635334 438566 635434
rect 438666 635334 438790 635434
rect 438890 635334 438924 635434
rect 437764 635210 438924 635334
rect 437764 635110 437894 635210
rect 437994 635110 438118 635210
rect 438218 635110 438342 635210
rect 438442 635110 438566 635210
rect 438666 635110 438790 635210
rect 438890 635110 438924 635210
rect 437764 634986 438924 635110
rect 437764 634886 437894 634986
rect 437994 634886 438118 634986
rect 438218 634886 438342 634986
rect 438442 634886 438566 634986
rect 438666 634886 438790 634986
rect 438890 634886 438924 634986
rect 437764 634762 438924 634886
rect 437764 634662 437894 634762
rect 437994 634662 438118 634762
rect 438218 634662 438342 634762
rect 438442 634662 438566 634762
rect 438666 634662 438790 634762
rect 438890 634662 438924 634762
rect 437764 634538 438924 634662
rect 437764 634438 437894 634538
rect 437994 634438 438118 634538
rect 438218 634438 438342 634538
rect 438442 634438 438566 634538
rect 438666 634438 438790 634538
rect 438890 634438 438924 634538
rect 437764 634314 438924 634438
rect 437764 634214 437894 634314
rect 437994 634214 438118 634314
rect 438218 634214 438342 634314
rect 438442 634214 438566 634314
rect 438666 634214 438790 634314
rect 438890 634214 438924 634314
rect 437764 634090 438924 634214
rect 437764 633990 437894 634090
rect 437994 633990 438118 634090
rect 438218 633990 438342 634090
rect 438442 633990 438566 634090
rect 438666 633990 438790 634090
rect 438890 633990 438924 634090
rect 437764 633866 438924 633990
rect 437764 633766 437894 633866
rect 437994 633766 438118 633866
rect 438218 633766 438342 633866
rect 438442 633766 438566 633866
rect 438666 633766 438790 633866
rect 438890 633766 438924 633866
rect 437764 633642 438924 633766
rect 437764 633542 437894 633642
rect 437994 633542 438118 633642
rect 438218 633542 438342 633642
rect 438442 633542 438566 633642
rect 438666 633542 438790 633642
rect 438890 633542 438924 633642
rect 437764 633418 438924 633542
rect 437764 633318 437894 633418
rect 437994 633318 438118 633418
rect 438218 633318 438342 633418
rect 438442 633318 438566 633418
rect 438666 633318 438790 633418
rect 438890 633318 438924 633418
rect 437764 633194 438924 633318
rect 437764 633094 437894 633194
rect 437994 633094 438118 633194
rect 438218 633094 438342 633194
rect 438442 633094 438566 633194
rect 438666 633094 438790 633194
rect 438890 633094 438924 633194
rect 437764 632970 438924 633094
rect 437764 632870 437894 632970
rect 437994 632870 438118 632970
rect 438218 632870 438342 632970
rect 438442 632870 438566 632970
rect 438666 632870 438790 632970
rect 438890 632870 438924 632970
rect 437764 632746 438924 632870
rect 437764 632646 437894 632746
rect 437994 632646 438118 632746
rect 438218 632646 438342 632746
rect 438442 632646 438566 632746
rect 438666 632646 438790 632746
rect 438890 632646 438924 632746
rect 437764 632522 438924 632646
rect 437764 632422 437894 632522
rect 437994 632422 438118 632522
rect 438218 632422 438342 632522
rect 438442 632422 438566 632522
rect 438666 632422 438790 632522
rect 438890 632422 438924 632522
rect 437764 632298 438924 632422
rect 437764 632198 437894 632298
rect 437994 632198 438118 632298
rect 438218 632198 438342 632298
rect 438442 632198 438566 632298
rect 438666 632198 438790 632298
rect 438890 632198 438924 632298
rect 437764 632074 438924 632198
rect 437764 631974 437894 632074
rect 437994 631974 438118 632074
rect 438218 631974 438342 632074
rect 438442 631974 438566 632074
rect 438666 631974 438790 632074
rect 438890 631974 438924 632074
rect 443628 632331 444268 632337
rect 443628 632051 443634 632331
rect 444262 632051 444268 632331
rect 443628 632045 444268 632051
rect 437764 631850 438924 631974
rect 437764 631750 437894 631850
rect 437994 631750 438118 631850
rect 438218 631750 438342 631850
rect 438442 631750 438566 631850
rect 438666 631750 438790 631850
rect 438890 631750 438924 631850
rect 437764 631626 438924 631750
rect 437764 631526 437894 631626
rect 437994 631526 438118 631626
rect 438218 631526 438342 631626
rect 438442 631526 438566 631626
rect 438666 631526 438790 631626
rect 438890 631526 438924 631626
rect 437764 631402 438924 631526
rect 437764 631302 437894 631402
rect 437994 631302 438118 631402
rect 438218 631302 438342 631402
rect 438442 631302 438566 631402
rect 438666 631302 438790 631402
rect 438890 631302 438924 631402
rect 437764 631178 438924 631302
rect 437764 631078 437894 631178
rect 437994 631078 438118 631178
rect 438218 631078 438342 631178
rect 438442 631078 438566 631178
rect 438666 631078 438790 631178
rect 438890 631078 438924 631178
rect 437764 630954 438924 631078
rect 437764 630854 437894 630954
rect 437994 630854 438118 630954
rect 438218 630854 438342 630954
rect 438442 630854 438566 630954
rect 438666 630854 438790 630954
rect 438890 630854 438924 630954
rect 437764 630730 438924 630854
rect 437764 630630 437894 630730
rect 437994 630630 438118 630730
rect 438218 630630 438342 630730
rect 438442 630630 438566 630730
rect 438666 630630 438790 630730
rect 438890 630630 438924 630730
rect 437764 630506 438924 630630
rect 437764 630406 437894 630506
rect 437994 630406 438118 630506
rect 438218 630406 438342 630506
rect 438442 630406 438566 630506
rect 438666 630406 438790 630506
rect 438890 630406 438924 630506
rect 437764 630282 438924 630406
rect 437764 630182 437894 630282
rect 437994 630182 438118 630282
rect 438218 630182 438342 630282
rect 438442 630182 438566 630282
rect 438666 630182 438790 630282
rect 438890 630182 438924 630282
rect 437764 630126 438924 630182
rect 444360 629250 451530 637482
rect 482144 636782 483230 636788
rect 482044 636778 483230 636782
rect 482044 636678 482174 636778
rect 482274 636678 482398 636778
rect 482498 636678 482622 636778
rect 482722 636678 482846 636778
rect 482946 636678 483070 636778
rect 483170 636678 483230 636778
rect 482044 636554 483230 636678
rect 482044 636454 482174 636554
rect 482274 636454 482398 636554
rect 482498 636454 482622 636554
rect 482722 636454 482846 636554
rect 482946 636454 483070 636554
rect 483170 636454 483230 636554
rect 482044 636330 483230 636454
rect 482044 636230 482174 636330
rect 482274 636230 482398 636330
rect 482498 636230 482622 636330
rect 482722 636230 482846 636330
rect 482946 636230 483070 636330
rect 483170 636230 483230 636330
rect 482044 636106 483230 636230
rect 482044 636006 482174 636106
rect 482274 636006 482398 636106
rect 482498 636006 482622 636106
rect 482722 636006 482846 636106
rect 482946 636006 483070 636106
rect 483170 636006 483230 636106
rect 482044 635882 483230 636006
rect 482044 635782 482174 635882
rect 482274 635782 482398 635882
rect 482498 635782 482622 635882
rect 482722 635782 482846 635882
rect 482946 635782 483070 635882
rect 483170 635782 483230 635882
rect 482044 635658 483230 635782
rect 482044 635558 482174 635658
rect 482274 635558 482398 635658
rect 482498 635558 482622 635658
rect 482722 635558 482846 635658
rect 482946 635558 483070 635658
rect 483170 635558 483230 635658
rect 482044 635434 483230 635558
rect 482044 635334 482174 635434
rect 482274 635334 482398 635434
rect 482498 635334 482622 635434
rect 482722 635334 482846 635434
rect 482946 635334 483070 635434
rect 483170 635334 483230 635434
rect 482044 635210 483230 635334
rect 482044 635110 482174 635210
rect 482274 635110 482398 635210
rect 482498 635110 482622 635210
rect 482722 635110 482846 635210
rect 482946 635110 483070 635210
rect 483170 635110 483230 635210
rect 482044 634986 483230 635110
rect 482044 634886 482174 634986
rect 482274 634886 482398 634986
rect 482498 634886 482622 634986
rect 482722 634886 482846 634986
rect 482946 634886 483070 634986
rect 483170 634886 483230 634986
rect 482044 634762 483230 634886
rect 482044 634662 482174 634762
rect 482274 634662 482398 634762
rect 482498 634662 482622 634762
rect 482722 634662 482846 634762
rect 482946 634662 483070 634762
rect 483170 634662 483230 634762
rect 482044 634538 483230 634662
rect 482044 634438 482174 634538
rect 482274 634438 482398 634538
rect 482498 634438 482622 634538
rect 482722 634438 482846 634538
rect 482946 634438 483070 634538
rect 483170 634438 483230 634538
rect 482044 634314 483230 634438
rect 482044 634214 482174 634314
rect 482274 634214 482398 634314
rect 482498 634214 482622 634314
rect 482722 634214 482846 634314
rect 482946 634214 483070 634314
rect 483170 634214 483230 634314
rect 482044 634090 483230 634214
rect 482044 633990 482174 634090
rect 482274 633990 482398 634090
rect 482498 633990 482622 634090
rect 482722 633990 482846 634090
rect 482946 633990 483070 634090
rect 483170 633990 483230 634090
rect 482044 633866 483230 633990
rect 482044 633766 482174 633866
rect 482274 633766 482398 633866
rect 482498 633766 482622 633866
rect 482722 633766 482846 633866
rect 482946 633766 483070 633866
rect 483170 633766 483230 633866
rect 482044 633642 483230 633766
rect 482044 633542 482174 633642
rect 482274 633542 482398 633642
rect 482498 633542 482622 633642
rect 482722 633542 482846 633642
rect 482946 633542 483070 633642
rect 483170 633542 483230 633642
rect 482044 633418 483230 633542
rect 482044 633318 482174 633418
rect 482274 633318 482398 633418
rect 482498 633318 482622 633418
rect 482722 633318 482846 633418
rect 482946 633318 483070 633418
rect 483170 633318 483230 633418
rect 482044 633194 483230 633318
rect 482044 633094 482174 633194
rect 482274 633094 482398 633194
rect 482498 633094 482622 633194
rect 482722 633094 482846 633194
rect 482946 633094 483070 633194
rect 483170 633094 483230 633194
rect 482044 632970 483230 633094
rect 482044 632870 482174 632970
rect 482274 632870 482398 632970
rect 482498 632870 482622 632970
rect 482722 632870 482846 632970
rect 482946 632870 483070 632970
rect 483170 632870 483230 632970
rect 482044 632746 483230 632870
rect 482044 632646 482174 632746
rect 482274 632646 482398 632746
rect 482498 632646 482622 632746
rect 482722 632646 482846 632746
rect 482946 632646 483070 632746
rect 483170 632646 483230 632746
rect 482044 632522 483230 632646
rect 482044 632422 482174 632522
rect 482274 632422 482398 632522
rect 482498 632422 482622 632522
rect 482722 632422 482846 632522
rect 482946 632422 483070 632522
rect 483170 632422 483230 632522
rect 452119 632331 452759 632337
rect 452119 632051 452125 632331
rect 452753 632051 452759 632331
rect 452119 632045 452759 632051
rect 482044 632298 483230 632422
rect 482044 632198 482174 632298
rect 482274 632198 482398 632298
rect 482498 632198 482622 632298
rect 482722 632198 482846 632298
rect 482946 632198 483070 632298
rect 483170 632198 483230 632298
rect 482044 632074 483230 632198
rect 482044 631974 482174 632074
rect 482274 631974 482398 632074
rect 482498 631974 482622 632074
rect 482722 631974 482846 632074
rect 482946 631974 483070 632074
rect 483170 631974 483230 632074
rect 482044 631850 483230 631974
rect 482044 631750 482174 631850
rect 482274 631750 482398 631850
rect 482498 631750 482622 631850
rect 482722 631750 482846 631850
rect 482946 631750 483070 631850
rect 483170 631750 483230 631850
rect 482044 631626 483230 631750
rect 482044 631526 482174 631626
rect 482274 631526 482398 631626
rect 482498 631526 482622 631626
rect 482722 631526 482846 631626
rect 482946 631526 483070 631626
rect 483170 631526 483230 631626
rect 482044 631402 483230 631526
rect 482044 631302 482174 631402
rect 482274 631302 482398 631402
rect 482498 631302 482622 631402
rect 482722 631302 482846 631402
rect 482946 631302 483070 631402
rect 483170 631302 483230 631402
rect 482044 631178 483230 631302
rect 482044 631078 482174 631178
rect 482274 631078 482398 631178
rect 482498 631078 482622 631178
rect 482722 631078 482846 631178
rect 482946 631078 483070 631178
rect 483170 631078 483230 631178
rect 482044 630954 483230 631078
rect 482044 630854 482174 630954
rect 482274 630854 482398 630954
rect 482498 630854 482622 630954
rect 482722 630854 482846 630954
rect 482946 630854 483070 630954
rect 483170 630854 483230 630954
rect 482044 630730 483230 630854
rect 482044 630630 482174 630730
rect 482274 630630 482398 630730
rect 482498 630630 482622 630730
rect 482722 630630 482846 630730
rect 482946 630630 483070 630730
rect 483170 630630 483230 630730
rect 482044 630506 483230 630630
rect 482044 630406 482174 630506
rect 482274 630406 482398 630506
rect 482498 630406 482622 630506
rect 482722 630406 482846 630506
rect 482946 630406 483070 630506
rect 483170 630406 483230 630506
rect 482044 630282 483230 630406
rect 482044 630182 482174 630282
rect 482274 630182 482398 630282
rect 482498 630182 482622 630282
rect 482722 630182 482846 630282
rect 482946 630182 483070 630282
rect 483170 630182 483230 630282
rect 482044 630126 483230 630182
rect 486272 636344 492928 644000
rect 486272 630600 487200 636344
rect 491984 630600 492928 636344
rect 442982 629244 470713 629250
rect 442982 629130 442990 629244
rect 452236 629130 470713 629244
rect 441982 629028 470713 629130
rect 441982 629022 470714 629028
rect 441982 629012 470724 629022
rect 441982 628694 452754 629012
rect 470692 628694 470724 629012
rect 441982 628688 470724 628694
rect 444360 628654 451530 628688
rect 428964 617202 429964 622946
rect 434748 617202 435620 622946
rect 428964 616702 435620 617202
rect 438864 627656 456004 627702
rect 438864 627556 438920 627656
rect 439020 627556 439144 627656
rect 439244 627556 439368 627656
rect 439468 627556 439592 627656
rect 439692 627556 439816 627656
rect 439916 627556 440040 627656
rect 440140 627556 440264 627656
rect 440364 627556 440488 627656
rect 440588 627556 440712 627656
rect 440812 627556 440936 627656
rect 441036 627556 441160 627656
rect 441260 627556 441384 627656
rect 441484 627556 441608 627656
rect 441708 627556 441832 627656
rect 441932 627556 442056 627656
rect 442156 627556 442280 627656
rect 442380 627556 442504 627656
rect 442604 627556 442728 627656
rect 442828 627556 442952 627656
rect 443052 627556 443176 627656
rect 443276 627556 443400 627656
rect 443500 627556 443624 627656
rect 443724 627556 443848 627656
rect 443948 627556 444072 627656
rect 444172 627556 444296 627656
rect 444396 627556 444520 627656
rect 444620 627556 444744 627656
rect 444844 627556 444968 627656
rect 445068 627556 445192 627656
rect 445292 627556 445416 627656
rect 445516 627556 449390 627656
rect 449490 627556 449614 627656
rect 449714 627556 449838 627656
rect 449938 627556 450062 627656
rect 450162 627556 450286 627656
rect 450386 627556 450510 627656
rect 450610 627556 450734 627656
rect 450834 627556 450958 627656
rect 451058 627556 451182 627656
rect 451282 627556 451406 627656
rect 451506 627556 451630 627656
rect 451730 627556 451854 627656
rect 451954 627556 452078 627656
rect 452178 627556 452302 627656
rect 452402 627556 452526 627656
rect 452626 627556 452750 627656
rect 452850 627556 452974 627656
rect 453074 627556 453198 627656
rect 453298 627556 453422 627656
rect 453522 627556 453646 627656
rect 453746 627556 453870 627656
rect 453970 627556 454094 627656
rect 454194 627556 454318 627656
rect 454418 627556 454542 627656
rect 454642 627556 454766 627656
rect 454866 627556 454990 627656
rect 455090 627556 455214 627656
rect 455314 627556 455438 627656
rect 455538 627556 455662 627656
rect 455762 627556 455886 627656
rect 455986 627556 456004 627656
rect 438864 627432 456004 627556
rect 438864 627332 438920 627432
rect 439020 627332 439144 627432
rect 439244 627332 439368 627432
rect 439468 627332 439592 627432
rect 439692 627332 439816 627432
rect 439916 627332 440040 627432
rect 440140 627332 440264 627432
rect 440364 627332 440488 627432
rect 440588 627332 440712 627432
rect 440812 627332 440936 627432
rect 441036 627332 441160 627432
rect 441260 627332 441384 627432
rect 441484 627332 441608 627432
rect 441708 627332 441832 627432
rect 441932 627332 442056 627432
rect 442156 627332 442280 627432
rect 442380 627332 442504 627432
rect 442604 627332 442728 627432
rect 442828 627332 442952 627432
rect 443052 627332 443176 627432
rect 443276 627332 443400 627432
rect 443500 627332 443624 627432
rect 443724 627332 443848 627432
rect 443948 627332 444072 627432
rect 444172 627332 444296 627432
rect 444396 627332 444520 627432
rect 444620 627332 444744 627432
rect 444844 627332 444968 627432
rect 445068 627332 445192 627432
rect 445292 627332 445416 627432
rect 445516 627332 449390 627432
rect 449490 627332 449614 627432
rect 449714 627332 449838 627432
rect 449938 627332 450062 627432
rect 450162 627332 450286 627432
rect 450386 627332 450510 627432
rect 450610 627332 450734 627432
rect 450834 627332 450958 627432
rect 451058 627332 451182 627432
rect 451282 627332 451406 627432
rect 451506 627332 451630 627432
rect 451730 627332 451854 627432
rect 451954 627332 452078 627432
rect 452178 627332 452302 627432
rect 452402 627332 452526 627432
rect 452626 627332 452750 627432
rect 452850 627332 452974 627432
rect 453074 627332 453198 627432
rect 453298 627332 453422 627432
rect 453522 627332 453646 627432
rect 453746 627332 453870 627432
rect 453970 627332 454094 627432
rect 454194 627332 454318 627432
rect 454418 627332 454542 627432
rect 454642 627332 454766 627432
rect 454866 627332 454990 627432
rect 455090 627332 455214 627432
rect 455314 627332 455438 627432
rect 455538 627332 455662 627432
rect 455762 627332 455886 627432
rect 455986 627332 456004 627432
rect 438864 627208 456004 627332
rect 438864 627108 438920 627208
rect 439020 627108 439144 627208
rect 439244 627108 439368 627208
rect 439468 627108 439592 627208
rect 439692 627108 439816 627208
rect 439916 627108 440040 627208
rect 440140 627108 440264 627208
rect 440364 627108 440488 627208
rect 440588 627108 440712 627208
rect 440812 627108 440936 627208
rect 441036 627108 441160 627208
rect 441260 627108 441384 627208
rect 441484 627108 441608 627208
rect 441708 627108 441832 627208
rect 441932 627108 442056 627208
rect 442156 627108 442280 627208
rect 442380 627108 442504 627208
rect 442604 627108 442728 627208
rect 442828 627108 442952 627208
rect 443052 627108 443176 627208
rect 443276 627108 443400 627208
rect 443500 627108 443624 627208
rect 443724 627108 443848 627208
rect 443948 627108 444072 627208
rect 444172 627108 444296 627208
rect 444396 627108 444520 627208
rect 444620 627108 444744 627208
rect 444844 627108 444968 627208
rect 445068 627108 445192 627208
rect 445292 627108 445416 627208
rect 445516 627108 449390 627208
rect 449490 627108 449614 627208
rect 449714 627108 449838 627208
rect 449938 627108 450062 627208
rect 450162 627108 450286 627208
rect 450386 627108 450510 627208
rect 450610 627108 450734 627208
rect 450834 627108 450958 627208
rect 451058 627108 451182 627208
rect 451282 627108 451406 627208
rect 451506 627108 451630 627208
rect 451730 627108 451854 627208
rect 451954 627108 452078 627208
rect 452178 627108 452302 627208
rect 452402 627108 452526 627208
rect 452626 627108 452750 627208
rect 452850 627108 452974 627208
rect 453074 627108 453198 627208
rect 453298 627108 453422 627208
rect 453522 627108 453646 627208
rect 453746 627108 453870 627208
rect 453970 627108 454094 627208
rect 454194 627108 454318 627208
rect 454418 627108 454542 627208
rect 454642 627108 454766 627208
rect 454866 627108 454990 627208
rect 455090 627108 455214 627208
rect 455314 627108 455438 627208
rect 455538 627108 455662 627208
rect 455762 627108 455886 627208
rect 455986 627108 456004 627208
rect 438864 626984 456004 627108
rect 438864 626884 438920 626984
rect 439020 626884 439144 626984
rect 439244 626884 439368 626984
rect 439468 626884 439592 626984
rect 439692 626884 439816 626984
rect 439916 626884 440040 626984
rect 440140 626884 440264 626984
rect 440364 626884 440488 626984
rect 440588 626884 440712 626984
rect 440812 626884 440936 626984
rect 441036 626884 441160 626984
rect 441260 626884 441384 626984
rect 441484 626884 441608 626984
rect 441708 626884 441832 626984
rect 441932 626884 442056 626984
rect 442156 626884 442280 626984
rect 442380 626884 442504 626984
rect 442604 626884 442728 626984
rect 442828 626884 442952 626984
rect 443052 626884 443176 626984
rect 443276 626884 443400 626984
rect 443500 626884 443624 626984
rect 443724 626884 443848 626984
rect 443948 626884 444072 626984
rect 444172 626884 444296 626984
rect 444396 626884 444520 626984
rect 444620 626884 444744 626984
rect 444844 626884 444968 626984
rect 445068 626884 445192 626984
rect 445292 626884 445416 626984
rect 445516 626884 449390 626984
rect 449490 626884 449614 626984
rect 449714 626884 449838 626984
rect 449938 626884 450062 626984
rect 450162 626884 450286 626984
rect 450386 626884 450510 626984
rect 450610 626884 450734 626984
rect 450834 626884 450958 626984
rect 451058 626884 451182 626984
rect 451282 626884 451406 626984
rect 451506 626884 451630 626984
rect 451730 626884 451854 626984
rect 451954 626884 452078 626984
rect 452178 626884 452302 626984
rect 452402 626884 452526 626984
rect 452626 626884 452750 626984
rect 452850 626884 452974 626984
rect 453074 626884 453198 626984
rect 453298 626884 453422 626984
rect 453522 626884 453646 626984
rect 453746 626884 453870 626984
rect 453970 626884 454094 626984
rect 454194 626884 454318 626984
rect 454418 626884 454542 626984
rect 454642 626884 454766 626984
rect 454866 626884 454990 626984
rect 455090 626884 455214 626984
rect 455314 626884 455438 626984
rect 455538 626884 455662 626984
rect 455762 626884 455886 626984
rect 455986 626884 456004 626984
rect 438864 626760 456004 626884
rect 438864 626660 438920 626760
rect 439020 626660 439144 626760
rect 439244 626660 439368 626760
rect 439468 626660 439592 626760
rect 439692 626660 439816 626760
rect 439916 626660 440040 626760
rect 440140 626660 440264 626760
rect 440364 626660 440488 626760
rect 440588 626660 440712 626760
rect 440812 626660 440936 626760
rect 441036 626660 441160 626760
rect 441260 626660 441384 626760
rect 441484 626660 441608 626760
rect 441708 626660 441832 626760
rect 441932 626660 442056 626760
rect 442156 626660 442280 626760
rect 442380 626660 442504 626760
rect 442604 626660 442728 626760
rect 442828 626660 442952 626760
rect 443052 626660 443176 626760
rect 443276 626660 443400 626760
rect 443500 626660 443624 626760
rect 443724 626660 443848 626760
rect 443948 626660 444072 626760
rect 444172 626660 444296 626760
rect 444396 626660 444520 626760
rect 444620 626660 444744 626760
rect 444844 626660 444968 626760
rect 445068 626660 445192 626760
rect 445292 626660 445416 626760
rect 445516 626660 449390 626760
rect 449490 626660 449614 626760
rect 449714 626660 449838 626760
rect 449938 626660 450062 626760
rect 450162 626660 450286 626760
rect 450386 626660 450510 626760
rect 450610 626660 450734 626760
rect 450834 626660 450958 626760
rect 451058 626660 451182 626760
rect 451282 626660 451406 626760
rect 451506 626660 451630 626760
rect 451730 626660 451854 626760
rect 451954 626660 452078 626760
rect 452178 626660 452302 626760
rect 452402 626660 452526 626760
rect 452626 626660 452750 626760
rect 452850 626660 452974 626760
rect 453074 626660 453198 626760
rect 453298 626660 453422 626760
rect 453522 626660 453646 626760
rect 453746 626660 453870 626760
rect 453970 626660 454094 626760
rect 454194 626660 454318 626760
rect 454418 626660 454542 626760
rect 454642 626660 454766 626760
rect 454866 626660 454990 626760
rect 455090 626660 455214 626760
rect 455314 626660 455438 626760
rect 455538 626660 455662 626760
rect 455762 626660 455886 626760
rect 455986 626660 456004 626760
rect 438864 625282 456004 626660
rect 438864 623262 456024 625282
rect 438864 617518 438964 623262
rect 443748 617518 444964 623262
rect 449748 617518 450964 623262
rect 455748 617518 456024 623262
rect 438864 616702 456024 617518
rect 457004 609506 470724 628688
rect 475604 627676 482444 627722
rect 475604 627576 475660 627676
rect 475760 627576 475884 627676
rect 475984 627576 476108 627676
rect 476208 627576 476332 627676
rect 476432 627576 476556 627676
rect 476656 627576 476780 627676
rect 476880 627576 477004 627676
rect 477104 627576 477228 627676
rect 477328 627576 477452 627676
rect 477552 627576 477676 627676
rect 477776 627576 477900 627676
rect 478000 627576 478124 627676
rect 478224 627576 478348 627676
rect 478448 627576 478572 627676
rect 478672 627576 478796 627676
rect 478896 627576 479020 627676
rect 479120 627576 479244 627676
rect 479344 627576 479468 627676
rect 479568 627576 479692 627676
rect 479792 627576 479916 627676
rect 480016 627576 480140 627676
rect 480240 627576 480364 627676
rect 480464 627576 480588 627676
rect 480688 627576 480812 627676
rect 480912 627576 481036 627676
rect 481136 627576 481260 627676
rect 481360 627576 481484 627676
rect 481584 627576 481708 627676
rect 481808 627576 481932 627676
rect 482032 627576 482156 627676
rect 482256 627576 482444 627676
rect 475604 627452 482444 627576
rect 475604 627352 475660 627452
rect 475760 627352 475884 627452
rect 475984 627352 476108 627452
rect 476208 627352 476332 627452
rect 476432 627352 476556 627452
rect 476656 627352 476780 627452
rect 476880 627352 477004 627452
rect 477104 627352 477228 627452
rect 477328 627352 477452 627452
rect 477552 627352 477676 627452
rect 477776 627352 477900 627452
rect 478000 627352 478124 627452
rect 478224 627352 478348 627452
rect 478448 627352 478572 627452
rect 478672 627352 478796 627452
rect 478896 627352 479020 627452
rect 479120 627352 479244 627452
rect 479344 627352 479468 627452
rect 479568 627352 479692 627452
rect 479792 627352 479916 627452
rect 480016 627352 480140 627452
rect 480240 627352 480364 627452
rect 480464 627352 480588 627452
rect 480688 627352 480812 627452
rect 480912 627352 481036 627452
rect 481136 627352 481260 627452
rect 481360 627352 481484 627452
rect 481584 627352 481708 627452
rect 481808 627352 481932 627452
rect 482032 627352 482156 627452
rect 482256 627352 482444 627452
rect 475604 627228 482444 627352
rect 475604 627128 475660 627228
rect 475760 627128 475884 627228
rect 475984 627128 476108 627228
rect 476208 627128 476332 627228
rect 476432 627128 476556 627228
rect 476656 627128 476780 627228
rect 476880 627128 477004 627228
rect 477104 627128 477228 627228
rect 477328 627128 477452 627228
rect 477552 627128 477676 627228
rect 477776 627128 477900 627228
rect 478000 627128 478124 627228
rect 478224 627128 478348 627228
rect 478448 627128 478572 627228
rect 478672 627128 478796 627228
rect 478896 627128 479020 627228
rect 479120 627128 479244 627228
rect 479344 627128 479468 627228
rect 479568 627128 479692 627228
rect 479792 627128 479916 627228
rect 480016 627128 480140 627228
rect 480240 627128 480364 627228
rect 480464 627128 480588 627228
rect 480688 627128 480812 627228
rect 480912 627128 481036 627228
rect 481136 627128 481260 627228
rect 481360 627128 481484 627228
rect 481584 627128 481708 627228
rect 481808 627128 481932 627228
rect 482032 627128 482156 627228
rect 482256 627128 482444 627228
rect 475604 627004 482444 627128
rect 475604 626904 475660 627004
rect 475760 626904 475884 627004
rect 475984 626904 476108 627004
rect 476208 626904 476332 627004
rect 476432 626904 476556 627004
rect 476656 626904 476780 627004
rect 476880 626904 477004 627004
rect 477104 626904 477228 627004
rect 477328 626904 477452 627004
rect 477552 626904 477676 627004
rect 477776 626904 477900 627004
rect 478000 626904 478124 627004
rect 478224 626904 478348 627004
rect 478448 626904 478572 627004
rect 478672 626904 478796 627004
rect 478896 626904 479020 627004
rect 479120 626904 479244 627004
rect 479344 626904 479468 627004
rect 479568 626904 479692 627004
rect 479792 626904 479916 627004
rect 480016 626904 480140 627004
rect 480240 626904 480364 627004
rect 480464 626904 480588 627004
rect 480688 626904 480812 627004
rect 480912 626904 481036 627004
rect 481136 626904 481260 627004
rect 481360 626904 481484 627004
rect 481584 626904 481708 627004
rect 481808 626904 481932 627004
rect 482032 626904 482156 627004
rect 482256 626904 482444 627004
rect 475604 626780 482444 626904
rect 475604 626680 475660 626780
rect 475760 626680 475884 626780
rect 475984 626680 476108 626780
rect 476208 626680 476332 626780
rect 476432 626680 476556 626780
rect 476656 626680 476780 626780
rect 476880 626680 477004 626780
rect 477104 626680 477228 626780
rect 477328 626680 477452 626780
rect 477552 626680 477676 626780
rect 477776 626680 477900 626780
rect 478000 626680 478124 626780
rect 478224 626680 478348 626780
rect 478448 626680 478572 626780
rect 478672 626680 478796 626780
rect 478896 626680 479020 626780
rect 479120 626680 479244 626780
rect 479344 626680 479468 626780
rect 479568 626680 479692 626780
rect 479792 626680 479916 626780
rect 480016 626680 480140 626780
rect 480240 626680 480364 626780
rect 480464 626680 480588 626780
rect 480688 626680 480812 626780
rect 480912 626680 481036 626780
rect 481136 626680 481260 626780
rect 481360 626680 481484 626780
rect 481584 626680 481708 626780
rect 481808 626680 481932 626780
rect 482032 626680 482156 626780
rect 482256 626680 482444 626780
rect 475604 626646 482444 626680
rect 475624 623266 482444 626646
rect 475624 617522 476524 623266
rect 481308 617522 482444 623266
rect 475624 616902 482444 617522
rect 486272 623144 492928 630600
rect 486272 617400 487200 623144
rect 491984 617400 492928 623144
rect 486272 616744 492928 617400
rect 457004 603762 457524 609506
rect 462308 603762 465524 609506
rect 470308 603762 470724 609506
rect 457004 603262 470724 603762
<< via3 >>
rect 429964 657022 434748 662766
rect 438964 657022 443748 662766
rect 444964 657022 449748 662766
rect 450964 657022 455748 662766
rect 438920 654776 439020 654876
rect 439144 654776 439244 654876
rect 439368 654776 439468 654876
rect 439592 654776 439692 654876
rect 439816 654776 439916 654876
rect 440040 654776 440140 654876
rect 440264 654776 440364 654876
rect 440488 654776 440588 654876
rect 440712 654776 440812 654876
rect 440936 654776 441036 654876
rect 441160 654776 441260 654876
rect 441384 654776 441484 654876
rect 441608 654776 441708 654876
rect 441832 654776 441932 654876
rect 442056 654776 442156 654876
rect 442280 654776 442380 654876
rect 442504 654776 442604 654876
rect 442728 654776 442828 654876
rect 442952 654776 443052 654876
rect 443176 654776 443276 654876
rect 443400 654776 443500 654876
rect 443624 654776 443724 654876
rect 443848 654776 443948 654876
rect 444072 654776 444172 654876
rect 444296 654776 444396 654876
rect 444520 654776 444620 654876
rect 444744 654776 444844 654876
rect 444968 654776 445068 654876
rect 445192 654776 445292 654876
rect 445416 654776 445516 654876
rect 449390 654776 449490 654876
rect 449614 654776 449714 654876
rect 449838 654776 449938 654876
rect 450062 654776 450162 654876
rect 450286 654776 450386 654876
rect 450510 654776 450610 654876
rect 450734 654776 450834 654876
rect 450958 654776 451058 654876
rect 451182 654776 451282 654876
rect 451406 654776 451506 654876
rect 451630 654776 451730 654876
rect 451854 654776 451954 654876
rect 452078 654776 452178 654876
rect 452302 654776 452402 654876
rect 452526 654776 452626 654876
rect 452750 654776 452850 654876
rect 452974 654776 453074 654876
rect 453198 654776 453298 654876
rect 453422 654776 453522 654876
rect 453646 654776 453746 654876
rect 453870 654776 453970 654876
rect 454094 654776 454194 654876
rect 454318 654776 454418 654876
rect 454542 654776 454642 654876
rect 454766 654776 454866 654876
rect 454990 654776 455090 654876
rect 455214 654776 455314 654876
rect 455438 654776 455538 654876
rect 455662 654776 455762 654876
rect 455886 654776 455986 654876
rect 438920 654552 439020 654652
rect 439144 654552 439244 654652
rect 439368 654552 439468 654652
rect 439592 654552 439692 654652
rect 439816 654552 439916 654652
rect 440040 654552 440140 654652
rect 440264 654552 440364 654652
rect 440488 654552 440588 654652
rect 440712 654552 440812 654652
rect 440936 654552 441036 654652
rect 441160 654552 441260 654652
rect 441384 654552 441484 654652
rect 441608 654552 441708 654652
rect 441832 654552 441932 654652
rect 442056 654552 442156 654652
rect 442280 654552 442380 654652
rect 442504 654552 442604 654652
rect 442728 654552 442828 654652
rect 442952 654552 443052 654652
rect 443176 654552 443276 654652
rect 443400 654552 443500 654652
rect 443624 654552 443724 654652
rect 443848 654552 443948 654652
rect 444072 654552 444172 654652
rect 444296 654552 444396 654652
rect 444520 654552 444620 654652
rect 444744 654552 444844 654652
rect 444968 654552 445068 654652
rect 445192 654552 445292 654652
rect 445416 654552 445516 654652
rect 449390 654552 449490 654652
rect 449614 654552 449714 654652
rect 449838 654552 449938 654652
rect 450062 654552 450162 654652
rect 450286 654552 450386 654652
rect 450510 654552 450610 654652
rect 450734 654552 450834 654652
rect 450958 654552 451058 654652
rect 451182 654552 451282 654652
rect 451406 654552 451506 654652
rect 451630 654552 451730 654652
rect 451854 654552 451954 654652
rect 452078 654552 452178 654652
rect 452302 654552 452402 654652
rect 452526 654552 452626 654652
rect 452750 654552 452850 654652
rect 452974 654552 453074 654652
rect 453198 654552 453298 654652
rect 453422 654552 453522 654652
rect 453646 654552 453746 654652
rect 453870 654552 453970 654652
rect 454094 654552 454194 654652
rect 454318 654552 454418 654652
rect 454542 654552 454642 654652
rect 454766 654552 454866 654652
rect 454990 654552 455090 654652
rect 455214 654552 455314 654652
rect 455438 654552 455538 654652
rect 455662 654552 455762 654652
rect 455886 654552 455986 654652
rect 438920 654328 439020 654428
rect 439144 654328 439244 654428
rect 439368 654328 439468 654428
rect 439592 654328 439692 654428
rect 439816 654328 439916 654428
rect 440040 654328 440140 654428
rect 440264 654328 440364 654428
rect 440488 654328 440588 654428
rect 440712 654328 440812 654428
rect 440936 654328 441036 654428
rect 441160 654328 441260 654428
rect 441384 654328 441484 654428
rect 441608 654328 441708 654428
rect 441832 654328 441932 654428
rect 442056 654328 442156 654428
rect 442280 654328 442380 654428
rect 442504 654328 442604 654428
rect 442728 654328 442828 654428
rect 442952 654328 443052 654428
rect 443176 654328 443276 654428
rect 443400 654328 443500 654428
rect 443624 654328 443724 654428
rect 443848 654328 443948 654428
rect 444072 654328 444172 654428
rect 444296 654328 444396 654428
rect 444520 654328 444620 654428
rect 444744 654328 444844 654428
rect 444968 654328 445068 654428
rect 445192 654328 445292 654428
rect 445416 654328 445516 654428
rect 449390 654328 449490 654428
rect 449614 654328 449714 654428
rect 449838 654328 449938 654428
rect 450062 654328 450162 654428
rect 450286 654328 450386 654428
rect 450510 654328 450610 654428
rect 450734 654328 450834 654428
rect 450958 654328 451058 654428
rect 451182 654328 451282 654428
rect 451406 654328 451506 654428
rect 451630 654328 451730 654428
rect 451854 654328 451954 654428
rect 452078 654328 452178 654428
rect 452302 654328 452402 654428
rect 452526 654328 452626 654428
rect 452750 654328 452850 654428
rect 452974 654328 453074 654428
rect 453198 654328 453298 654428
rect 453422 654328 453522 654428
rect 453646 654328 453746 654428
rect 453870 654328 453970 654428
rect 454094 654328 454194 654428
rect 454318 654328 454418 654428
rect 454542 654328 454642 654428
rect 454766 654328 454866 654428
rect 454990 654328 455090 654428
rect 455214 654328 455314 654428
rect 455438 654328 455538 654428
rect 455662 654328 455762 654428
rect 455886 654328 455986 654428
rect 438920 654104 439020 654204
rect 439144 654104 439244 654204
rect 439368 654104 439468 654204
rect 439592 654104 439692 654204
rect 439816 654104 439916 654204
rect 440040 654104 440140 654204
rect 440264 654104 440364 654204
rect 440488 654104 440588 654204
rect 440712 654104 440812 654204
rect 440936 654104 441036 654204
rect 441160 654104 441260 654204
rect 441384 654104 441484 654204
rect 441608 654104 441708 654204
rect 441832 654104 441932 654204
rect 442056 654104 442156 654204
rect 442280 654104 442380 654204
rect 442504 654104 442604 654204
rect 442728 654104 442828 654204
rect 442952 654104 443052 654204
rect 443176 654104 443276 654204
rect 443400 654104 443500 654204
rect 443624 654104 443724 654204
rect 443848 654104 443948 654204
rect 444072 654104 444172 654204
rect 444296 654104 444396 654204
rect 444520 654104 444620 654204
rect 444744 654104 444844 654204
rect 444968 654104 445068 654204
rect 445192 654104 445292 654204
rect 445416 654104 445516 654204
rect 449390 654104 449490 654204
rect 449614 654104 449714 654204
rect 449838 654104 449938 654204
rect 450062 654104 450162 654204
rect 450286 654104 450386 654204
rect 450510 654104 450610 654204
rect 450734 654104 450834 654204
rect 450958 654104 451058 654204
rect 451182 654104 451282 654204
rect 451406 654104 451506 654204
rect 451630 654104 451730 654204
rect 451854 654104 451954 654204
rect 452078 654104 452178 654204
rect 452302 654104 452402 654204
rect 452526 654104 452626 654204
rect 452750 654104 452850 654204
rect 452974 654104 453074 654204
rect 453198 654104 453298 654204
rect 453422 654104 453522 654204
rect 453646 654104 453746 654204
rect 453870 654104 453970 654204
rect 454094 654104 454194 654204
rect 454318 654104 454418 654204
rect 454542 654104 454642 654204
rect 454766 654104 454866 654204
rect 454990 654104 455090 654204
rect 455214 654104 455314 654204
rect 455438 654104 455538 654204
rect 455662 654104 455762 654204
rect 455886 654104 455986 654204
rect 438920 653880 439020 653980
rect 439144 653880 439244 653980
rect 439368 653880 439468 653980
rect 439592 653880 439692 653980
rect 439816 653880 439916 653980
rect 440040 653880 440140 653980
rect 440264 653880 440364 653980
rect 440488 653880 440588 653980
rect 440712 653880 440812 653980
rect 440936 653880 441036 653980
rect 441160 653880 441260 653980
rect 441384 653880 441484 653980
rect 441608 653880 441708 653980
rect 441832 653880 441932 653980
rect 442056 653880 442156 653980
rect 442280 653880 442380 653980
rect 442504 653880 442604 653980
rect 442728 653880 442828 653980
rect 442952 653880 443052 653980
rect 443176 653880 443276 653980
rect 443400 653880 443500 653980
rect 443624 653880 443724 653980
rect 443848 653880 443948 653980
rect 444072 653880 444172 653980
rect 444296 653880 444396 653980
rect 444520 653880 444620 653980
rect 444744 653880 444844 653980
rect 444968 653880 445068 653980
rect 445192 653880 445292 653980
rect 445416 653880 445516 653980
rect 449390 653880 449490 653980
rect 449614 653880 449714 653980
rect 449838 653880 449938 653980
rect 450062 653880 450162 653980
rect 450286 653880 450386 653980
rect 450510 653880 450610 653980
rect 450734 653880 450834 653980
rect 450958 653880 451058 653980
rect 451182 653880 451282 653980
rect 451406 653880 451506 653980
rect 451630 653880 451730 653980
rect 451854 653880 451954 653980
rect 452078 653880 452178 653980
rect 452302 653880 452402 653980
rect 452526 653880 452626 653980
rect 452750 653880 452850 653980
rect 452974 653880 453074 653980
rect 453198 653880 453298 653980
rect 453422 653880 453522 653980
rect 453646 653880 453746 653980
rect 453870 653880 453970 653980
rect 454094 653880 454194 653980
rect 454318 653880 454418 653980
rect 454542 653880 454642 653980
rect 454766 653880 454866 653980
rect 454990 653880 455090 653980
rect 455214 653880 455314 653980
rect 455438 653880 455538 653980
rect 455662 653880 455762 653980
rect 455886 653880 455986 653980
rect 440687 652760 451961 652769
rect 440687 651922 440696 652760
rect 440696 651922 451952 652760
rect 451952 651922 451961 652760
rect 440687 651913 451961 651922
rect 429964 643622 434748 649366
rect 437894 650078 437994 650178
rect 438118 650078 438218 650178
rect 438342 650078 438442 650178
rect 438566 650078 438666 650178
rect 438790 650078 438890 650178
rect 437894 649854 437994 649954
rect 438118 649854 438218 649954
rect 438342 649854 438442 649954
rect 438566 649854 438666 649954
rect 438790 649854 438890 649954
rect 437894 649630 437994 649730
rect 438118 649630 438218 649730
rect 438342 649630 438442 649730
rect 438566 649630 438666 649730
rect 438790 649630 438890 649730
rect 437894 649406 437994 649506
rect 438118 649406 438218 649506
rect 438342 649406 438442 649506
rect 438566 649406 438666 649506
rect 438790 649406 438890 649506
rect 437894 649182 437994 649282
rect 438118 649182 438218 649282
rect 438342 649182 438442 649282
rect 438566 649182 438666 649282
rect 438790 649182 438890 649282
rect 437894 648958 437994 649058
rect 438118 648958 438218 649058
rect 438342 648958 438442 649058
rect 438566 648958 438666 649058
rect 438790 648958 438890 649058
rect 437894 648734 437994 648834
rect 438118 648734 438218 648834
rect 438342 648734 438442 648834
rect 438566 648734 438666 648834
rect 438790 648734 438890 648834
rect 437894 648510 437994 648610
rect 438118 648510 438218 648610
rect 438342 648510 438442 648610
rect 438566 648510 438666 648610
rect 438790 648510 438890 648610
rect 437894 648286 437994 648386
rect 438118 648286 438218 648386
rect 438342 648286 438442 648386
rect 438566 648286 438666 648386
rect 438790 648286 438890 648386
rect 437894 648062 437994 648162
rect 438118 648062 438218 648162
rect 438342 648062 438442 648162
rect 438566 648062 438666 648162
rect 438790 648062 438890 648162
rect 437894 647838 437994 647938
rect 438118 647838 438218 647938
rect 438342 647838 438442 647938
rect 438566 647838 438666 647938
rect 438790 647838 438890 647938
rect 437894 647614 437994 647714
rect 438118 647614 438218 647714
rect 438342 647614 438442 647714
rect 438566 647614 438666 647714
rect 438790 647614 438890 647714
rect 437894 647390 437994 647490
rect 438118 647390 438218 647490
rect 438342 647390 438442 647490
rect 438566 647390 438666 647490
rect 438790 647390 438890 647490
rect 437894 647166 437994 647266
rect 438118 647166 438218 647266
rect 438342 647166 438442 647266
rect 438566 647166 438666 647266
rect 438790 647166 438890 647266
rect 437894 646942 437994 647042
rect 438118 646942 438218 647042
rect 438342 646942 438442 647042
rect 438566 646942 438666 647042
rect 438790 646942 438890 647042
rect 437894 646718 437994 646818
rect 438118 646718 438218 646818
rect 438342 646718 438442 646818
rect 438566 646718 438666 646818
rect 438790 646718 438890 646818
rect 437894 646494 437994 646594
rect 438118 646494 438218 646594
rect 438342 646494 438442 646594
rect 438566 646494 438666 646594
rect 438790 646494 438890 646594
rect 437894 646270 437994 646370
rect 438118 646270 438218 646370
rect 438342 646270 438442 646370
rect 438566 646270 438666 646370
rect 438790 646270 438890 646370
rect 437894 646046 437994 646146
rect 438118 646046 438218 646146
rect 438342 646046 438442 646146
rect 438566 646046 438666 646146
rect 438790 646046 438890 646146
rect 437894 645822 437994 645922
rect 438118 645822 438218 645922
rect 438342 645822 438442 645922
rect 438566 645822 438666 645922
rect 438790 645822 438890 645922
rect 437894 645598 437994 645698
rect 438118 645598 438218 645698
rect 438342 645598 438442 645698
rect 438566 645598 438666 645698
rect 438790 645598 438890 645698
rect 437894 645374 437994 645474
rect 438118 645374 438218 645474
rect 438342 645374 438442 645474
rect 438566 645374 438666 645474
rect 438790 645374 438890 645474
rect 437894 645150 437994 645250
rect 438118 645150 438218 645250
rect 438342 645150 438442 645250
rect 438566 645150 438666 645250
rect 438790 645150 438890 645250
rect 437894 644926 437994 645026
rect 438118 644926 438218 645026
rect 438342 644926 438442 645026
rect 438566 644926 438666 645026
rect 438790 644926 438890 645026
rect 437894 644702 437994 644802
rect 438118 644702 438218 644802
rect 438342 644702 438442 644802
rect 438566 644702 438666 644802
rect 438790 644702 438890 644802
rect 437894 644478 437994 644578
rect 438118 644478 438218 644578
rect 438342 644478 438442 644578
rect 438566 644478 438666 644578
rect 438790 644478 438890 644578
rect 437894 644254 437994 644354
rect 438118 644254 438218 644354
rect 438342 644254 438442 644354
rect 438566 644254 438666 644354
rect 438790 644254 438890 644354
rect 437894 644030 437994 644130
rect 438118 644030 438218 644130
rect 438342 644030 438442 644130
rect 438566 644030 438666 644130
rect 438790 644030 438890 644130
rect 437894 643806 437994 643906
rect 438118 643806 438218 643906
rect 438342 643806 438442 643906
rect 438566 643806 438666 643906
rect 438790 643806 438890 643906
rect 437894 643582 437994 643682
rect 438118 643582 438218 643682
rect 438342 643582 438442 643682
rect 438566 643582 438666 643682
rect 438790 643582 438890 643682
rect 444975 643782 445039 644326
rect 445694 643782 445758 644326
rect 446413 643782 446477 644326
rect 447132 643782 447196 644326
rect 447851 643782 447915 644326
rect 448570 643782 448634 644326
rect 449289 643782 449353 644326
rect 450008 643782 450072 644326
rect 450727 643782 450791 644326
rect 451446 643782 451510 644326
rect 444975 643082 445039 643626
rect 445694 643082 445758 643626
rect 446413 643082 446477 643626
rect 447132 643082 447196 643626
rect 447851 643082 447915 643626
rect 448570 643082 448634 643626
rect 449289 643082 449353 643626
rect 450008 643082 450072 643626
rect 450727 643082 450791 643626
rect 451446 643082 451510 643626
rect 444975 642382 445039 642926
rect 445694 642382 445758 642926
rect 446413 642382 446477 642926
rect 447132 642382 447196 642926
rect 447851 642382 447915 642926
rect 448570 642382 448634 642926
rect 449289 642382 449353 642926
rect 450008 642382 450072 642926
rect 450727 642382 450791 642926
rect 451446 642382 451510 642926
rect 444975 641682 445039 642226
rect 445694 641682 445758 642226
rect 446413 641682 446477 642226
rect 447132 641682 447196 642226
rect 447851 641682 447915 642226
rect 448570 641682 448634 642226
rect 449289 641682 449353 642226
rect 450008 641682 450072 642226
rect 450727 641682 450791 642226
rect 451446 641682 451510 642226
rect 444975 640982 445039 641526
rect 445694 640982 445758 641526
rect 446413 640982 446477 641526
rect 447132 640982 447196 641526
rect 447851 640982 447915 641526
rect 448570 640982 448634 641526
rect 449289 640982 449353 641526
rect 450008 640982 450072 641526
rect 450727 640982 450791 641526
rect 451446 640982 451510 641526
rect 444975 640282 445039 640826
rect 445694 640282 445758 640826
rect 446413 640282 446477 640826
rect 447132 640282 447196 640826
rect 447851 640282 447915 640826
rect 448570 640282 448634 640826
rect 449289 640282 449353 640826
rect 450008 640282 450072 640826
rect 450727 640282 450791 640826
rect 451446 640282 451510 640826
rect 444975 639582 445039 640126
rect 445694 639582 445758 640126
rect 446413 639582 446477 640126
rect 447132 639582 447196 640126
rect 447851 639582 447915 640126
rect 448570 639582 448634 640126
rect 449289 639582 449353 640126
rect 450008 639582 450072 640126
rect 450727 639582 450791 640126
rect 451446 639582 451510 640126
rect 476524 657342 481308 663086
rect 475660 654796 475760 654896
rect 475884 654796 475984 654896
rect 476108 654796 476208 654896
rect 476332 654796 476432 654896
rect 476556 654796 476656 654896
rect 476780 654796 476880 654896
rect 477004 654796 477104 654896
rect 477228 654796 477328 654896
rect 477452 654796 477552 654896
rect 477676 654796 477776 654896
rect 477900 654796 478000 654896
rect 478124 654796 478224 654896
rect 478348 654796 478448 654896
rect 478572 654796 478672 654896
rect 478796 654796 478896 654896
rect 479020 654796 479120 654896
rect 479244 654796 479344 654896
rect 479468 654796 479568 654896
rect 479692 654796 479792 654896
rect 479916 654796 480016 654896
rect 480140 654796 480240 654896
rect 480364 654796 480464 654896
rect 480588 654796 480688 654896
rect 480812 654796 480912 654896
rect 481036 654796 481136 654896
rect 481260 654796 481360 654896
rect 481484 654796 481584 654896
rect 481708 654796 481808 654896
rect 481932 654796 482032 654896
rect 482156 654796 482256 654896
rect 475660 654572 475760 654672
rect 475884 654572 475984 654672
rect 476108 654572 476208 654672
rect 476332 654572 476432 654672
rect 476556 654572 476656 654672
rect 476780 654572 476880 654672
rect 477004 654572 477104 654672
rect 477228 654572 477328 654672
rect 477452 654572 477552 654672
rect 477676 654572 477776 654672
rect 477900 654572 478000 654672
rect 478124 654572 478224 654672
rect 478348 654572 478448 654672
rect 478572 654572 478672 654672
rect 478796 654572 478896 654672
rect 479020 654572 479120 654672
rect 479244 654572 479344 654672
rect 479468 654572 479568 654672
rect 479692 654572 479792 654672
rect 479916 654572 480016 654672
rect 480140 654572 480240 654672
rect 480364 654572 480464 654672
rect 480588 654572 480688 654672
rect 480812 654572 480912 654672
rect 481036 654572 481136 654672
rect 481260 654572 481360 654672
rect 481484 654572 481584 654672
rect 481708 654572 481808 654672
rect 481932 654572 482032 654672
rect 482156 654572 482256 654672
rect 475660 654348 475760 654448
rect 475884 654348 475984 654448
rect 476108 654348 476208 654448
rect 476332 654348 476432 654448
rect 476556 654348 476656 654448
rect 476780 654348 476880 654448
rect 477004 654348 477104 654448
rect 477228 654348 477328 654448
rect 477452 654348 477552 654448
rect 477676 654348 477776 654448
rect 477900 654348 478000 654448
rect 478124 654348 478224 654448
rect 478348 654348 478448 654448
rect 478572 654348 478672 654448
rect 478796 654348 478896 654448
rect 479020 654348 479120 654448
rect 479244 654348 479344 654448
rect 479468 654348 479568 654448
rect 479692 654348 479792 654448
rect 479916 654348 480016 654448
rect 480140 654348 480240 654448
rect 480364 654348 480464 654448
rect 480588 654348 480688 654448
rect 480812 654348 480912 654448
rect 481036 654348 481136 654448
rect 481260 654348 481360 654448
rect 481484 654348 481584 654448
rect 481708 654348 481808 654448
rect 481932 654348 482032 654448
rect 482156 654348 482256 654448
rect 475660 654124 475760 654224
rect 475884 654124 475984 654224
rect 476108 654124 476208 654224
rect 476332 654124 476432 654224
rect 476556 654124 476656 654224
rect 476780 654124 476880 654224
rect 477004 654124 477104 654224
rect 477228 654124 477328 654224
rect 477452 654124 477552 654224
rect 477676 654124 477776 654224
rect 477900 654124 478000 654224
rect 478124 654124 478224 654224
rect 478348 654124 478448 654224
rect 478572 654124 478672 654224
rect 478796 654124 478896 654224
rect 479020 654124 479120 654224
rect 479244 654124 479344 654224
rect 479468 654124 479568 654224
rect 479692 654124 479792 654224
rect 479916 654124 480016 654224
rect 480140 654124 480240 654224
rect 480364 654124 480464 654224
rect 480588 654124 480688 654224
rect 480812 654124 480912 654224
rect 481036 654124 481136 654224
rect 481260 654124 481360 654224
rect 481484 654124 481584 654224
rect 481708 654124 481808 654224
rect 481932 654124 482032 654224
rect 482156 654124 482256 654224
rect 475660 653900 475760 654000
rect 475884 653900 475984 654000
rect 476108 653900 476208 654000
rect 476332 653900 476432 654000
rect 476556 653900 476656 654000
rect 476780 653900 476880 654000
rect 477004 653900 477104 654000
rect 477228 653900 477328 654000
rect 477452 653900 477552 654000
rect 477676 653900 477776 654000
rect 477900 653900 478000 654000
rect 478124 653900 478224 654000
rect 478348 653900 478448 654000
rect 478572 653900 478672 654000
rect 478796 653900 478896 654000
rect 479020 653900 479120 654000
rect 479244 653900 479344 654000
rect 479468 653900 479568 654000
rect 479692 653900 479792 654000
rect 479916 653900 480016 654000
rect 480140 653900 480240 654000
rect 480364 653900 480464 654000
rect 480588 653900 480688 654000
rect 480812 653900 480912 654000
rect 481036 653900 481136 654000
rect 481260 653900 481360 654000
rect 481484 653900 481584 654000
rect 481708 653900 481808 654000
rect 481932 653900 482032 654000
rect 482156 653900 482256 654000
rect 487200 657400 491984 663144
rect 482174 650078 482274 650178
rect 482398 650078 482498 650178
rect 482622 650078 482722 650178
rect 482846 650078 482946 650178
rect 483070 650078 483170 650178
rect 482174 649854 482274 649954
rect 482398 649854 482498 649954
rect 482622 649854 482722 649954
rect 482846 649854 482946 649954
rect 483070 649854 483170 649954
rect 482174 649630 482274 649730
rect 482398 649630 482498 649730
rect 482622 649630 482722 649730
rect 482846 649630 482946 649730
rect 483070 649630 483170 649730
rect 482174 649406 482274 649506
rect 482398 649406 482498 649506
rect 482622 649406 482722 649506
rect 482846 649406 482946 649506
rect 483070 649406 483170 649506
rect 482174 649182 482274 649282
rect 482398 649182 482498 649282
rect 482622 649182 482722 649282
rect 482846 649182 482946 649282
rect 483070 649182 483170 649282
rect 482174 648958 482274 649058
rect 482398 648958 482498 649058
rect 482622 648958 482722 649058
rect 482846 648958 482946 649058
rect 483070 648958 483170 649058
rect 482174 648734 482274 648834
rect 482398 648734 482498 648834
rect 482622 648734 482722 648834
rect 482846 648734 482946 648834
rect 483070 648734 483170 648834
rect 482174 648510 482274 648610
rect 482398 648510 482498 648610
rect 482622 648510 482722 648610
rect 482846 648510 482946 648610
rect 483070 648510 483170 648610
rect 482174 648286 482274 648386
rect 482398 648286 482498 648386
rect 482622 648286 482722 648386
rect 482846 648286 482946 648386
rect 483070 648286 483170 648386
rect 482174 648062 482274 648162
rect 482398 648062 482498 648162
rect 482622 648062 482722 648162
rect 482846 648062 482946 648162
rect 483070 648062 483170 648162
rect 482174 647838 482274 647938
rect 482398 647838 482498 647938
rect 482622 647838 482722 647938
rect 482846 647838 482946 647938
rect 483070 647838 483170 647938
rect 482174 647614 482274 647714
rect 482398 647614 482498 647714
rect 482622 647614 482722 647714
rect 482846 647614 482946 647714
rect 483070 647614 483170 647714
rect 482174 647390 482274 647490
rect 482398 647390 482498 647490
rect 482622 647390 482722 647490
rect 482846 647390 482946 647490
rect 483070 647390 483170 647490
rect 482174 647166 482274 647266
rect 482398 647166 482498 647266
rect 482622 647166 482722 647266
rect 482846 647166 482946 647266
rect 483070 647166 483170 647266
rect 482174 646942 482274 647042
rect 482398 646942 482498 647042
rect 482622 646942 482722 647042
rect 482846 646942 482946 647042
rect 483070 646942 483170 647042
rect 482174 646718 482274 646818
rect 482398 646718 482498 646818
rect 482622 646718 482722 646818
rect 482846 646718 482946 646818
rect 483070 646718 483170 646818
rect 482174 646494 482274 646594
rect 482398 646494 482498 646594
rect 482622 646494 482722 646594
rect 482846 646494 482946 646594
rect 483070 646494 483170 646594
rect 482174 646270 482274 646370
rect 482398 646270 482498 646370
rect 482622 646270 482722 646370
rect 482846 646270 482946 646370
rect 483070 646270 483170 646370
rect 482174 646046 482274 646146
rect 482398 646046 482498 646146
rect 482622 646046 482722 646146
rect 482846 646046 482946 646146
rect 483070 646046 483170 646146
rect 482174 645822 482274 645922
rect 482398 645822 482498 645922
rect 482622 645822 482722 645922
rect 482846 645822 482946 645922
rect 483070 645822 483170 645922
rect 482174 645598 482274 645698
rect 482398 645598 482498 645698
rect 482622 645598 482722 645698
rect 482846 645598 482946 645698
rect 483070 645598 483170 645698
rect 482174 645374 482274 645474
rect 482398 645374 482498 645474
rect 482622 645374 482722 645474
rect 482846 645374 482946 645474
rect 483070 645374 483170 645474
rect 482174 645150 482274 645250
rect 482398 645150 482498 645250
rect 482622 645150 482722 645250
rect 482846 645150 482946 645250
rect 483070 645150 483170 645250
rect 482174 644926 482274 645026
rect 482398 644926 482498 645026
rect 482622 644926 482722 645026
rect 482846 644926 482946 645026
rect 483070 644926 483170 645026
rect 482174 644702 482274 644802
rect 482398 644702 482498 644802
rect 482622 644702 482722 644802
rect 482846 644702 482946 644802
rect 483070 644702 483170 644802
rect 482174 644478 482274 644578
rect 482398 644478 482498 644578
rect 482622 644478 482722 644578
rect 482846 644478 482946 644578
rect 483070 644478 483170 644578
rect 482174 644254 482274 644354
rect 482398 644254 482498 644354
rect 482622 644254 482722 644354
rect 482846 644254 482946 644354
rect 483070 644254 483170 644354
rect 482174 644030 482274 644130
rect 482398 644030 482498 644130
rect 482622 644030 482722 644130
rect 482846 644030 482946 644130
rect 483070 644030 483170 644130
rect 482174 643806 482274 643906
rect 482398 643806 482498 643906
rect 482622 643806 482722 643906
rect 482846 643806 482946 643906
rect 483070 643806 483170 643906
rect 482174 643582 482274 643682
rect 482398 643582 482498 643682
rect 482622 643582 482722 643682
rect 482846 643582 482946 643682
rect 483070 643582 483170 643682
rect 487200 644000 491984 649744
rect 459444 640850 459644 641050
rect 459878 640850 460078 641050
rect 460312 640850 460512 641050
rect 460746 640850 460946 641050
rect 461180 640850 461380 641050
rect 461614 640850 461814 641050
rect 462048 640850 462248 641050
rect 462482 640850 462682 641050
rect 462916 640850 463116 641050
rect 463350 640850 463550 641050
rect 463784 640850 463984 641050
rect 464184 640850 464384 641050
rect 464584 640850 464784 641050
rect 464984 640850 465184 641050
rect 465384 640850 465584 641050
rect 465784 640850 465984 641050
rect 466184 640850 466384 641050
rect 466584 640850 466784 641050
rect 466984 640850 467184 641050
rect 467384 640850 467584 641050
rect 468984 640850 469184 641050
rect 469384 640850 469584 641050
rect 469784 640850 469984 641050
rect 470184 640850 470384 641050
rect 470584 640850 470784 641050
rect 470984 640850 471184 641050
rect 471384 640850 471584 641050
rect 471784 640850 471984 641050
rect 472184 640850 472384 641050
rect 459444 640416 459644 640616
rect 459878 640416 460078 640616
rect 460312 640416 460512 640616
rect 460746 640416 460946 640616
rect 461180 640416 461380 640616
rect 461614 640416 461814 640616
rect 462048 640416 462248 640616
rect 462482 640416 462682 640616
rect 462916 640416 463116 640616
rect 463350 640416 463550 640616
rect 463784 640416 463984 640616
rect 459444 639982 459644 640182
rect 459878 639982 460078 640182
rect 460312 639982 460512 640182
rect 460746 639982 460946 640182
rect 461180 639982 461380 640182
rect 461614 639982 461814 640182
rect 462048 639982 462248 640182
rect 462482 639982 462682 640182
rect 462916 639982 463116 640182
rect 463350 639982 463550 640182
rect 463784 639982 463984 640182
rect 444975 638882 445039 639426
rect 445694 638882 445758 639426
rect 446413 638882 446477 639426
rect 447132 638882 447196 639426
rect 447851 638882 447915 639426
rect 448570 638882 448634 639426
rect 449289 638882 449353 639426
rect 450008 638882 450072 639426
rect 450727 638882 450791 639426
rect 451446 638882 451510 639426
rect 437900 638294 437964 638358
rect 438028 638294 438092 638358
rect 438156 638294 438220 638358
rect 438284 638294 438348 638358
rect 438412 638294 438476 638358
rect 438540 638294 438604 638358
rect 438668 638294 438732 638358
rect 438796 638294 438860 638358
rect 438924 638294 438988 638358
rect 437900 638166 437964 638230
rect 438028 638166 438092 638230
rect 438156 638166 438220 638230
rect 438284 638166 438348 638230
rect 438412 638166 438476 638230
rect 438540 638166 438604 638230
rect 438668 638166 438732 638230
rect 438796 638166 438860 638230
rect 438924 638166 438988 638230
rect 437900 638038 437964 638102
rect 438028 638038 438092 638102
rect 438156 638038 438220 638102
rect 438284 638038 438348 638102
rect 438412 638038 438476 638102
rect 438540 638038 438604 638102
rect 438668 638038 438732 638102
rect 438796 638038 438860 638102
rect 438924 638038 438988 638102
rect 437900 637910 437964 637974
rect 438028 637910 438092 637974
rect 438156 637910 438220 637974
rect 438284 637910 438348 637974
rect 438412 637910 438476 637974
rect 438540 637910 438604 637974
rect 438668 637910 438732 637974
rect 438796 637910 438860 637974
rect 438924 637910 438988 637974
rect 444975 638182 445039 638726
rect 445694 638182 445758 638726
rect 446413 638182 446477 638726
rect 447132 638182 447196 638726
rect 447851 638182 447915 638726
rect 448570 638182 448634 638726
rect 449289 638182 449353 638726
rect 450008 638182 450072 638726
rect 450727 638182 450791 638726
rect 451446 638182 451510 638726
rect 453002 638496 473312 639468
rect 444975 637482 445039 638026
rect 445694 637482 445758 638026
rect 446413 637482 446477 638026
rect 447132 637482 447196 638026
rect 447851 637482 447915 638026
rect 448570 637482 448634 638026
rect 449289 637482 449353 638026
rect 450008 637482 450072 638026
rect 450727 637482 450791 638026
rect 451446 637482 451510 638026
rect 429964 630222 434748 635966
rect 437894 636678 437994 636778
rect 438118 636678 438218 636778
rect 438342 636678 438442 636778
rect 438566 636678 438666 636778
rect 438790 636678 438890 636778
rect 437894 636454 437994 636554
rect 438118 636454 438218 636554
rect 438342 636454 438442 636554
rect 438566 636454 438666 636554
rect 438790 636454 438890 636554
rect 437894 636230 437994 636330
rect 438118 636230 438218 636330
rect 438342 636230 438442 636330
rect 438566 636230 438666 636330
rect 438790 636230 438890 636330
rect 437894 636006 437994 636106
rect 438118 636006 438218 636106
rect 438342 636006 438442 636106
rect 438566 636006 438666 636106
rect 438790 636006 438890 636106
rect 437894 635782 437994 635882
rect 438118 635782 438218 635882
rect 438342 635782 438442 635882
rect 438566 635782 438666 635882
rect 438790 635782 438890 635882
rect 437894 635558 437994 635658
rect 438118 635558 438218 635658
rect 438342 635558 438442 635658
rect 438566 635558 438666 635658
rect 438790 635558 438890 635658
rect 437894 635334 437994 635434
rect 438118 635334 438218 635434
rect 438342 635334 438442 635434
rect 438566 635334 438666 635434
rect 438790 635334 438890 635434
rect 437894 635110 437994 635210
rect 438118 635110 438218 635210
rect 438342 635110 438442 635210
rect 438566 635110 438666 635210
rect 438790 635110 438890 635210
rect 437894 634886 437994 634986
rect 438118 634886 438218 634986
rect 438342 634886 438442 634986
rect 438566 634886 438666 634986
rect 438790 634886 438890 634986
rect 437894 634662 437994 634762
rect 438118 634662 438218 634762
rect 438342 634662 438442 634762
rect 438566 634662 438666 634762
rect 438790 634662 438890 634762
rect 437894 634438 437994 634538
rect 438118 634438 438218 634538
rect 438342 634438 438442 634538
rect 438566 634438 438666 634538
rect 438790 634438 438890 634538
rect 437894 634214 437994 634314
rect 438118 634214 438218 634314
rect 438342 634214 438442 634314
rect 438566 634214 438666 634314
rect 438790 634214 438890 634314
rect 437894 633990 437994 634090
rect 438118 633990 438218 634090
rect 438342 633990 438442 634090
rect 438566 633990 438666 634090
rect 438790 633990 438890 634090
rect 437894 633766 437994 633866
rect 438118 633766 438218 633866
rect 438342 633766 438442 633866
rect 438566 633766 438666 633866
rect 438790 633766 438890 633866
rect 437894 633542 437994 633642
rect 438118 633542 438218 633642
rect 438342 633542 438442 633642
rect 438566 633542 438666 633642
rect 438790 633542 438890 633642
rect 437894 633318 437994 633418
rect 438118 633318 438218 633418
rect 438342 633318 438442 633418
rect 438566 633318 438666 633418
rect 438790 633318 438890 633418
rect 437894 633094 437994 633194
rect 438118 633094 438218 633194
rect 438342 633094 438442 633194
rect 438566 633094 438666 633194
rect 438790 633094 438890 633194
rect 437894 632870 437994 632970
rect 438118 632870 438218 632970
rect 438342 632870 438442 632970
rect 438566 632870 438666 632970
rect 438790 632870 438890 632970
rect 437894 632646 437994 632746
rect 438118 632646 438218 632746
rect 438342 632646 438442 632746
rect 438566 632646 438666 632746
rect 438790 632646 438890 632746
rect 437894 632422 437994 632522
rect 438118 632422 438218 632522
rect 438342 632422 438442 632522
rect 438566 632422 438666 632522
rect 438790 632422 438890 632522
rect 437894 632198 437994 632298
rect 438118 632198 438218 632298
rect 438342 632198 438442 632298
rect 438566 632198 438666 632298
rect 438790 632198 438890 632298
rect 437894 631974 437994 632074
rect 438118 631974 438218 632074
rect 438342 631974 438442 632074
rect 438566 631974 438666 632074
rect 438790 631974 438890 632074
rect 443634 632317 444262 632331
rect 443634 632065 443648 632317
rect 443648 632065 444248 632317
rect 444248 632065 444262 632317
rect 443634 632051 444262 632065
rect 437894 631750 437994 631850
rect 438118 631750 438218 631850
rect 438342 631750 438442 631850
rect 438566 631750 438666 631850
rect 438790 631750 438890 631850
rect 437894 631526 437994 631626
rect 438118 631526 438218 631626
rect 438342 631526 438442 631626
rect 438566 631526 438666 631626
rect 438790 631526 438890 631626
rect 437894 631302 437994 631402
rect 438118 631302 438218 631402
rect 438342 631302 438442 631402
rect 438566 631302 438666 631402
rect 438790 631302 438890 631402
rect 437894 631078 437994 631178
rect 438118 631078 438218 631178
rect 438342 631078 438442 631178
rect 438566 631078 438666 631178
rect 438790 631078 438890 631178
rect 437894 630854 437994 630954
rect 438118 630854 438218 630954
rect 438342 630854 438442 630954
rect 438566 630854 438666 630954
rect 438790 630854 438890 630954
rect 437894 630630 437994 630730
rect 438118 630630 438218 630730
rect 438342 630630 438442 630730
rect 438566 630630 438666 630730
rect 438790 630630 438890 630730
rect 437894 630406 437994 630506
rect 438118 630406 438218 630506
rect 438342 630406 438442 630506
rect 438566 630406 438666 630506
rect 438790 630406 438890 630506
rect 437894 630182 437994 630282
rect 438118 630182 438218 630282
rect 438342 630182 438442 630282
rect 438566 630182 438666 630282
rect 438790 630182 438890 630282
rect 482174 636678 482274 636778
rect 482398 636678 482498 636778
rect 482622 636678 482722 636778
rect 482846 636678 482946 636778
rect 483070 636678 483170 636778
rect 482174 636454 482274 636554
rect 482398 636454 482498 636554
rect 482622 636454 482722 636554
rect 482846 636454 482946 636554
rect 483070 636454 483170 636554
rect 482174 636230 482274 636330
rect 482398 636230 482498 636330
rect 482622 636230 482722 636330
rect 482846 636230 482946 636330
rect 483070 636230 483170 636330
rect 482174 636006 482274 636106
rect 482398 636006 482498 636106
rect 482622 636006 482722 636106
rect 482846 636006 482946 636106
rect 483070 636006 483170 636106
rect 482174 635782 482274 635882
rect 482398 635782 482498 635882
rect 482622 635782 482722 635882
rect 482846 635782 482946 635882
rect 483070 635782 483170 635882
rect 482174 635558 482274 635658
rect 482398 635558 482498 635658
rect 482622 635558 482722 635658
rect 482846 635558 482946 635658
rect 483070 635558 483170 635658
rect 482174 635334 482274 635434
rect 482398 635334 482498 635434
rect 482622 635334 482722 635434
rect 482846 635334 482946 635434
rect 483070 635334 483170 635434
rect 482174 635110 482274 635210
rect 482398 635110 482498 635210
rect 482622 635110 482722 635210
rect 482846 635110 482946 635210
rect 483070 635110 483170 635210
rect 482174 634886 482274 634986
rect 482398 634886 482498 634986
rect 482622 634886 482722 634986
rect 482846 634886 482946 634986
rect 483070 634886 483170 634986
rect 482174 634662 482274 634762
rect 482398 634662 482498 634762
rect 482622 634662 482722 634762
rect 482846 634662 482946 634762
rect 483070 634662 483170 634762
rect 482174 634438 482274 634538
rect 482398 634438 482498 634538
rect 482622 634438 482722 634538
rect 482846 634438 482946 634538
rect 483070 634438 483170 634538
rect 482174 634214 482274 634314
rect 482398 634214 482498 634314
rect 482622 634214 482722 634314
rect 482846 634214 482946 634314
rect 483070 634214 483170 634314
rect 482174 633990 482274 634090
rect 482398 633990 482498 634090
rect 482622 633990 482722 634090
rect 482846 633990 482946 634090
rect 483070 633990 483170 634090
rect 482174 633766 482274 633866
rect 482398 633766 482498 633866
rect 482622 633766 482722 633866
rect 482846 633766 482946 633866
rect 483070 633766 483170 633866
rect 482174 633542 482274 633642
rect 482398 633542 482498 633642
rect 482622 633542 482722 633642
rect 482846 633542 482946 633642
rect 483070 633542 483170 633642
rect 482174 633318 482274 633418
rect 482398 633318 482498 633418
rect 482622 633318 482722 633418
rect 482846 633318 482946 633418
rect 483070 633318 483170 633418
rect 482174 633094 482274 633194
rect 482398 633094 482498 633194
rect 482622 633094 482722 633194
rect 482846 633094 482946 633194
rect 483070 633094 483170 633194
rect 482174 632870 482274 632970
rect 482398 632870 482498 632970
rect 482622 632870 482722 632970
rect 482846 632870 482946 632970
rect 483070 632870 483170 632970
rect 482174 632646 482274 632746
rect 482398 632646 482498 632746
rect 482622 632646 482722 632746
rect 482846 632646 482946 632746
rect 483070 632646 483170 632746
rect 482174 632422 482274 632522
rect 482398 632422 482498 632522
rect 482622 632422 482722 632522
rect 482846 632422 482946 632522
rect 483070 632422 483170 632522
rect 452125 632317 452753 632331
rect 452125 632065 452139 632317
rect 452139 632065 452739 632317
rect 452739 632065 452753 632317
rect 452125 632051 452753 632065
rect 482174 632198 482274 632298
rect 482398 632198 482498 632298
rect 482622 632198 482722 632298
rect 482846 632198 482946 632298
rect 483070 632198 483170 632298
rect 482174 631974 482274 632074
rect 482398 631974 482498 632074
rect 482622 631974 482722 632074
rect 482846 631974 482946 632074
rect 483070 631974 483170 632074
rect 482174 631750 482274 631850
rect 482398 631750 482498 631850
rect 482622 631750 482722 631850
rect 482846 631750 482946 631850
rect 483070 631750 483170 631850
rect 482174 631526 482274 631626
rect 482398 631526 482498 631626
rect 482622 631526 482722 631626
rect 482846 631526 482946 631626
rect 483070 631526 483170 631626
rect 482174 631302 482274 631402
rect 482398 631302 482498 631402
rect 482622 631302 482722 631402
rect 482846 631302 482946 631402
rect 483070 631302 483170 631402
rect 482174 631078 482274 631178
rect 482398 631078 482498 631178
rect 482622 631078 482722 631178
rect 482846 631078 482946 631178
rect 483070 631078 483170 631178
rect 482174 630854 482274 630954
rect 482398 630854 482498 630954
rect 482622 630854 482722 630954
rect 482846 630854 482946 630954
rect 483070 630854 483170 630954
rect 482174 630630 482274 630730
rect 482398 630630 482498 630730
rect 482622 630630 482722 630730
rect 482846 630630 482946 630730
rect 483070 630630 483170 630730
rect 482174 630406 482274 630506
rect 482398 630406 482498 630506
rect 482622 630406 482722 630506
rect 482846 630406 482946 630506
rect 483070 630406 483170 630506
rect 482174 630182 482274 630282
rect 482398 630182 482498 630282
rect 482622 630182 482722 630282
rect 482846 630182 482946 630282
rect 483070 630182 483170 630282
rect 487200 630600 491984 636344
rect 429964 617202 434748 622946
rect 438920 627556 439020 627656
rect 439144 627556 439244 627656
rect 439368 627556 439468 627656
rect 439592 627556 439692 627656
rect 439816 627556 439916 627656
rect 440040 627556 440140 627656
rect 440264 627556 440364 627656
rect 440488 627556 440588 627656
rect 440712 627556 440812 627656
rect 440936 627556 441036 627656
rect 441160 627556 441260 627656
rect 441384 627556 441484 627656
rect 441608 627556 441708 627656
rect 441832 627556 441932 627656
rect 442056 627556 442156 627656
rect 442280 627556 442380 627656
rect 442504 627556 442604 627656
rect 442728 627556 442828 627656
rect 442952 627556 443052 627656
rect 443176 627556 443276 627656
rect 443400 627556 443500 627656
rect 443624 627556 443724 627656
rect 443848 627556 443948 627656
rect 444072 627556 444172 627656
rect 444296 627556 444396 627656
rect 444520 627556 444620 627656
rect 444744 627556 444844 627656
rect 444968 627556 445068 627656
rect 445192 627556 445292 627656
rect 445416 627556 445516 627656
rect 449390 627556 449490 627656
rect 449614 627556 449714 627656
rect 449838 627556 449938 627656
rect 450062 627556 450162 627656
rect 450286 627556 450386 627656
rect 450510 627556 450610 627656
rect 450734 627556 450834 627656
rect 450958 627556 451058 627656
rect 451182 627556 451282 627656
rect 451406 627556 451506 627656
rect 451630 627556 451730 627656
rect 451854 627556 451954 627656
rect 452078 627556 452178 627656
rect 452302 627556 452402 627656
rect 452526 627556 452626 627656
rect 452750 627556 452850 627656
rect 452974 627556 453074 627656
rect 453198 627556 453298 627656
rect 453422 627556 453522 627656
rect 453646 627556 453746 627656
rect 453870 627556 453970 627656
rect 454094 627556 454194 627656
rect 454318 627556 454418 627656
rect 454542 627556 454642 627656
rect 454766 627556 454866 627656
rect 454990 627556 455090 627656
rect 455214 627556 455314 627656
rect 455438 627556 455538 627656
rect 455662 627556 455762 627656
rect 455886 627556 455986 627656
rect 438920 627332 439020 627432
rect 439144 627332 439244 627432
rect 439368 627332 439468 627432
rect 439592 627332 439692 627432
rect 439816 627332 439916 627432
rect 440040 627332 440140 627432
rect 440264 627332 440364 627432
rect 440488 627332 440588 627432
rect 440712 627332 440812 627432
rect 440936 627332 441036 627432
rect 441160 627332 441260 627432
rect 441384 627332 441484 627432
rect 441608 627332 441708 627432
rect 441832 627332 441932 627432
rect 442056 627332 442156 627432
rect 442280 627332 442380 627432
rect 442504 627332 442604 627432
rect 442728 627332 442828 627432
rect 442952 627332 443052 627432
rect 443176 627332 443276 627432
rect 443400 627332 443500 627432
rect 443624 627332 443724 627432
rect 443848 627332 443948 627432
rect 444072 627332 444172 627432
rect 444296 627332 444396 627432
rect 444520 627332 444620 627432
rect 444744 627332 444844 627432
rect 444968 627332 445068 627432
rect 445192 627332 445292 627432
rect 445416 627332 445516 627432
rect 449390 627332 449490 627432
rect 449614 627332 449714 627432
rect 449838 627332 449938 627432
rect 450062 627332 450162 627432
rect 450286 627332 450386 627432
rect 450510 627332 450610 627432
rect 450734 627332 450834 627432
rect 450958 627332 451058 627432
rect 451182 627332 451282 627432
rect 451406 627332 451506 627432
rect 451630 627332 451730 627432
rect 451854 627332 451954 627432
rect 452078 627332 452178 627432
rect 452302 627332 452402 627432
rect 452526 627332 452626 627432
rect 452750 627332 452850 627432
rect 452974 627332 453074 627432
rect 453198 627332 453298 627432
rect 453422 627332 453522 627432
rect 453646 627332 453746 627432
rect 453870 627332 453970 627432
rect 454094 627332 454194 627432
rect 454318 627332 454418 627432
rect 454542 627332 454642 627432
rect 454766 627332 454866 627432
rect 454990 627332 455090 627432
rect 455214 627332 455314 627432
rect 455438 627332 455538 627432
rect 455662 627332 455762 627432
rect 455886 627332 455986 627432
rect 438920 627108 439020 627208
rect 439144 627108 439244 627208
rect 439368 627108 439468 627208
rect 439592 627108 439692 627208
rect 439816 627108 439916 627208
rect 440040 627108 440140 627208
rect 440264 627108 440364 627208
rect 440488 627108 440588 627208
rect 440712 627108 440812 627208
rect 440936 627108 441036 627208
rect 441160 627108 441260 627208
rect 441384 627108 441484 627208
rect 441608 627108 441708 627208
rect 441832 627108 441932 627208
rect 442056 627108 442156 627208
rect 442280 627108 442380 627208
rect 442504 627108 442604 627208
rect 442728 627108 442828 627208
rect 442952 627108 443052 627208
rect 443176 627108 443276 627208
rect 443400 627108 443500 627208
rect 443624 627108 443724 627208
rect 443848 627108 443948 627208
rect 444072 627108 444172 627208
rect 444296 627108 444396 627208
rect 444520 627108 444620 627208
rect 444744 627108 444844 627208
rect 444968 627108 445068 627208
rect 445192 627108 445292 627208
rect 445416 627108 445516 627208
rect 449390 627108 449490 627208
rect 449614 627108 449714 627208
rect 449838 627108 449938 627208
rect 450062 627108 450162 627208
rect 450286 627108 450386 627208
rect 450510 627108 450610 627208
rect 450734 627108 450834 627208
rect 450958 627108 451058 627208
rect 451182 627108 451282 627208
rect 451406 627108 451506 627208
rect 451630 627108 451730 627208
rect 451854 627108 451954 627208
rect 452078 627108 452178 627208
rect 452302 627108 452402 627208
rect 452526 627108 452626 627208
rect 452750 627108 452850 627208
rect 452974 627108 453074 627208
rect 453198 627108 453298 627208
rect 453422 627108 453522 627208
rect 453646 627108 453746 627208
rect 453870 627108 453970 627208
rect 454094 627108 454194 627208
rect 454318 627108 454418 627208
rect 454542 627108 454642 627208
rect 454766 627108 454866 627208
rect 454990 627108 455090 627208
rect 455214 627108 455314 627208
rect 455438 627108 455538 627208
rect 455662 627108 455762 627208
rect 455886 627108 455986 627208
rect 438920 626884 439020 626984
rect 439144 626884 439244 626984
rect 439368 626884 439468 626984
rect 439592 626884 439692 626984
rect 439816 626884 439916 626984
rect 440040 626884 440140 626984
rect 440264 626884 440364 626984
rect 440488 626884 440588 626984
rect 440712 626884 440812 626984
rect 440936 626884 441036 626984
rect 441160 626884 441260 626984
rect 441384 626884 441484 626984
rect 441608 626884 441708 626984
rect 441832 626884 441932 626984
rect 442056 626884 442156 626984
rect 442280 626884 442380 626984
rect 442504 626884 442604 626984
rect 442728 626884 442828 626984
rect 442952 626884 443052 626984
rect 443176 626884 443276 626984
rect 443400 626884 443500 626984
rect 443624 626884 443724 626984
rect 443848 626884 443948 626984
rect 444072 626884 444172 626984
rect 444296 626884 444396 626984
rect 444520 626884 444620 626984
rect 444744 626884 444844 626984
rect 444968 626884 445068 626984
rect 445192 626884 445292 626984
rect 445416 626884 445516 626984
rect 449390 626884 449490 626984
rect 449614 626884 449714 626984
rect 449838 626884 449938 626984
rect 450062 626884 450162 626984
rect 450286 626884 450386 626984
rect 450510 626884 450610 626984
rect 450734 626884 450834 626984
rect 450958 626884 451058 626984
rect 451182 626884 451282 626984
rect 451406 626884 451506 626984
rect 451630 626884 451730 626984
rect 451854 626884 451954 626984
rect 452078 626884 452178 626984
rect 452302 626884 452402 626984
rect 452526 626884 452626 626984
rect 452750 626884 452850 626984
rect 452974 626884 453074 626984
rect 453198 626884 453298 626984
rect 453422 626884 453522 626984
rect 453646 626884 453746 626984
rect 453870 626884 453970 626984
rect 454094 626884 454194 626984
rect 454318 626884 454418 626984
rect 454542 626884 454642 626984
rect 454766 626884 454866 626984
rect 454990 626884 455090 626984
rect 455214 626884 455314 626984
rect 455438 626884 455538 626984
rect 455662 626884 455762 626984
rect 455886 626884 455986 626984
rect 438920 626660 439020 626760
rect 439144 626660 439244 626760
rect 439368 626660 439468 626760
rect 439592 626660 439692 626760
rect 439816 626660 439916 626760
rect 440040 626660 440140 626760
rect 440264 626660 440364 626760
rect 440488 626660 440588 626760
rect 440712 626660 440812 626760
rect 440936 626660 441036 626760
rect 441160 626660 441260 626760
rect 441384 626660 441484 626760
rect 441608 626660 441708 626760
rect 441832 626660 441932 626760
rect 442056 626660 442156 626760
rect 442280 626660 442380 626760
rect 442504 626660 442604 626760
rect 442728 626660 442828 626760
rect 442952 626660 443052 626760
rect 443176 626660 443276 626760
rect 443400 626660 443500 626760
rect 443624 626660 443724 626760
rect 443848 626660 443948 626760
rect 444072 626660 444172 626760
rect 444296 626660 444396 626760
rect 444520 626660 444620 626760
rect 444744 626660 444844 626760
rect 444968 626660 445068 626760
rect 445192 626660 445292 626760
rect 445416 626660 445516 626760
rect 449390 626660 449490 626760
rect 449614 626660 449714 626760
rect 449838 626660 449938 626760
rect 450062 626660 450162 626760
rect 450286 626660 450386 626760
rect 450510 626660 450610 626760
rect 450734 626660 450834 626760
rect 450958 626660 451058 626760
rect 451182 626660 451282 626760
rect 451406 626660 451506 626760
rect 451630 626660 451730 626760
rect 451854 626660 451954 626760
rect 452078 626660 452178 626760
rect 452302 626660 452402 626760
rect 452526 626660 452626 626760
rect 452750 626660 452850 626760
rect 452974 626660 453074 626760
rect 453198 626660 453298 626760
rect 453422 626660 453522 626760
rect 453646 626660 453746 626760
rect 453870 626660 453970 626760
rect 454094 626660 454194 626760
rect 454318 626660 454418 626760
rect 454542 626660 454642 626760
rect 454766 626660 454866 626760
rect 454990 626660 455090 626760
rect 455214 626660 455314 626760
rect 455438 626660 455538 626760
rect 455662 626660 455762 626760
rect 455886 626660 455986 626760
rect 438964 617518 443748 623262
rect 444964 617518 449748 623262
rect 450964 617518 455748 623262
rect 475660 627576 475760 627676
rect 475884 627576 475984 627676
rect 476108 627576 476208 627676
rect 476332 627576 476432 627676
rect 476556 627576 476656 627676
rect 476780 627576 476880 627676
rect 477004 627576 477104 627676
rect 477228 627576 477328 627676
rect 477452 627576 477552 627676
rect 477676 627576 477776 627676
rect 477900 627576 478000 627676
rect 478124 627576 478224 627676
rect 478348 627576 478448 627676
rect 478572 627576 478672 627676
rect 478796 627576 478896 627676
rect 479020 627576 479120 627676
rect 479244 627576 479344 627676
rect 479468 627576 479568 627676
rect 479692 627576 479792 627676
rect 479916 627576 480016 627676
rect 480140 627576 480240 627676
rect 480364 627576 480464 627676
rect 480588 627576 480688 627676
rect 480812 627576 480912 627676
rect 481036 627576 481136 627676
rect 481260 627576 481360 627676
rect 481484 627576 481584 627676
rect 481708 627576 481808 627676
rect 481932 627576 482032 627676
rect 482156 627576 482256 627676
rect 475660 627352 475760 627452
rect 475884 627352 475984 627452
rect 476108 627352 476208 627452
rect 476332 627352 476432 627452
rect 476556 627352 476656 627452
rect 476780 627352 476880 627452
rect 477004 627352 477104 627452
rect 477228 627352 477328 627452
rect 477452 627352 477552 627452
rect 477676 627352 477776 627452
rect 477900 627352 478000 627452
rect 478124 627352 478224 627452
rect 478348 627352 478448 627452
rect 478572 627352 478672 627452
rect 478796 627352 478896 627452
rect 479020 627352 479120 627452
rect 479244 627352 479344 627452
rect 479468 627352 479568 627452
rect 479692 627352 479792 627452
rect 479916 627352 480016 627452
rect 480140 627352 480240 627452
rect 480364 627352 480464 627452
rect 480588 627352 480688 627452
rect 480812 627352 480912 627452
rect 481036 627352 481136 627452
rect 481260 627352 481360 627452
rect 481484 627352 481584 627452
rect 481708 627352 481808 627452
rect 481932 627352 482032 627452
rect 482156 627352 482256 627452
rect 475660 627128 475760 627228
rect 475884 627128 475984 627228
rect 476108 627128 476208 627228
rect 476332 627128 476432 627228
rect 476556 627128 476656 627228
rect 476780 627128 476880 627228
rect 477004 627128 477104 627228
rect 477228 627128 477328 627228
rect 477452 627128 477552 627228
rect 477676 627128 477776 627228
rect 477900 627128 478000 627228
rect 478124 627128 478224 627228
rect 478348 627128 478448 627228
rect 478572 627128 478672 627228
rect 478796 627128 478896 627228
rect 479020 627128 479120 627228
rect 479244 627128 479344 627228
rect 479468 627128 479568 627228
rect 479692 627128 479792 627228
rect 479916 627128 480016 627228
rect 480140 627128 480240 627228
rect 480364 627128 480464 627228
rect 480588 627128 480688 627228
rect 480812 627128 480912 627228
rect 481036 627128 481136 627228
rect 481260 627128 481360 627228
rect 481484 627128 481584 627228
rect 481708 627128 481808 627228
rect 481932 627128 482032 627228
rect 482156 627128 482256 627228
rect 475660 626904 475760 627004
rect 475884 626904 475984 627004
rect 476108 626904 476208 627004
rect 476332 626904 476432 627004
rect 476556 626904 476656 627004
rect 476780 626904 476880 627004
rect 477004 626904 477104 627004
rect 477228 626904 477328 627004
rect 477452 626904 477552 627004
rect 477676 626904 477776 627004
rect 477900 626904 478000 627004
rect 478124 626904 478224 627004
rect 478348 626904 478448 627004
rect 478572 626904 478672 627004
rect 478796 626904 478896 627004
rect 479020 626904 479120 627004
rect 479244 626904 479344 627004
rect 479468 626904 479568 627004
rect 479692 626904 479792 627004
rect 479916 626904 480016 627004
rect 480140 626904 480240 627004
rect 480364 626904 480464 627004
rect 480588 626904 480688 627004
rect 480812 626904 480912 627004
rect 481036 626904 481136 627004
rect 481260 626904 481360 627004
rect 481484 626904 481584 627004
rect 481708 626904 481808 627004
rect 481932 626904 482032 627004
rect 482156 626904 482256 627004
rect 475660 626680 475760 626780
rect 475884 626680 475984 626780
rect 476108 626680 476208 626780
rect 476332 626680 476432 626780
rect 476556 626680 476656 626780
rect 476780 626680 476880 626780
rect 477004 626680 477104 626780
rect 477228 626680 477328 626780
rect 477452 626680 477552 626780
rect 477676 626680 477776 626780
rect 477900 626680 478000 626780
rect 478124 626680 478224 626780
rect 478348 626680 478448 626780
rect 478572 626680 478672 626780
rect 478796 626680 478896 626780
rect 479020 626680 479120 626780
rect 479244 626680 479344 626780
rect 479468 626680 479568 626780
rect 479692 626680 479792 626780
rect 479916 626680 480016 626780
rect 480140 626680 480240 626780
rect 480364 626680 480464 626780
rect 480588 626680 480688 626780
rect 480812 626680 480912 626780
rect 481036 626680 481136 626780
rect 481260 626680 481360 626780
rect 481484 626680 481584 626780
rect 481708 626680 481808 626780
rect 481932 626680 482032 626780
rect 482156 626680 482256 626780
rect 476524 617522 481308 623266
rect 487200 617400 491984 623144
rect 457524 603762 462308 609506
rect 465524 603762 470308 609506
<< mimcap >>
rect 444460 644214 444860 644254
rect 444460 643894 444500 644214
rect 444820 643894 444860 644214
rect 444460 643854 444860 643894
rect 445179 644214 445579 644254
rect 445179 643894 445219 644214
rect 445539 643894 445579 644214
rect 445179 643854 445579 643894
rect 445898 644214 446298 644254
rect 445898 643894 445938 644214
rect 446258 643894 446298 644214
rect 445898 643854 446298 643894
rect 446617 644214 447017 644254
rect 446617 643894 446657 644214
rect 446977 643894 447017 644214
rect 446617 643854 447017 643894
rect 447336 644214 447736 644254
rect 447336 643894 447376 644214
rect 447696 643894 447736 644214
rect 447336 643854 447736 643894
rect 448055 644214 448455 644254
rect 448055 643894 448095 644214
rect 448415 643894 448455 644214
rect 448055 643854 448455 643894
rect 448774 644214 449174 644254
rect 448774 643894 448814 644214
rect 449134 643894 449174 644214
rect 448774 643854 449174 643894
rect 449493 644214 449893 644254
rect 449493 643894 449533 644214
rect 449853 643894 449893 644214
rect 449493 643854 449893 643894
rect 450212 644214 450612 644254
rect 450212 643894 450252 644214
rect 450572 643894 450612 644214
rect 450212 643854 450612 643894
rect 450931 644214 451331 644254
rect 450931 643894 450971 644214
rect 451291 643894 451331 644214
rect 450931 643854 451331 643894
rect 444460 643514 444860 643554
rect 444460 643194 444500 643514
rect 444820 643194 444860 643514
rect 444460 643154 444860 643194
rect 445179 643514 445579 643554
rect 445179 643194 445219 643514
rect 445539 643194 445579 643514
rect 445179 643154 445579 643194
rect 445898 643514 446298 643554
rect 445898 643194 445938 643514
rect 446258 643194 446298 643514
rect 445898 643154 446298 643194
rect 446617 643514 447017 643554
rect 446617 643194 446657 643514
rect 446977 643194 447017 643514
rect 446617 643154 447017 643194
rect 447336 643514 447736 643554
rect 447336 643194 447376 643514
rect 447696 643194 447736 643514
rect 447336 643154 447736 643194
rect 448055 643514 448455 643554
rect 448055 643194 448095 643514
rect 448415 643194 448455 643514
rect 448055 643154 448455 643194
rect 448774 643514 449174 643554
rect 448774 643194 448814 643514
rect 449134 643194 449174 643514
rect 448774 643154 449174 643194
rect 449493 643514 449893 643554
rect 449493 643194 449533 643514
rect 449853 643194 449893 643514
rect 449493 643154 449893 643194
rect 450212 643514 450612 643554
rect 450212 643194 450252 643514
rect 450572 643194 450612 643514
rect 450212 643154 450612 643194
rect 450931 643514 451331 643554
rect 450931 643194 450971 643514
rect 451291 643194 451331 643514
rect 450931 643154 451331 643194
rect 444460 642814 444860 642854
rect 444460 642494 444500 642814
rect 444820 642494 444860 642814
rect 444460 642454 444860 642494
rect 445179 642814 445579 642854
rect 445179 642494 445219 642814
rect 445539 642494 445579 642814
rect 445179 642454 445579 642494
rect 445898 642814 446298 642854
rect 445898 642494 445938 642814
rect 446258 642494 446298 642814
rect 445898 642454 446298 642494
rect 446617 642814 447017 642854
rect 446617 642494 446657 642814
rect 446977 642494 447017 642814
rect 446617 642454 447017 642494
rect 447336 642814 447736 642854
rect 447336 642494 447376 642814
rect 447696 642494 447736 642814
rect 447336 642454 447736 642494
rect 448055 642814 448455 642854
rect 448055 642494 448095 642814
rect 448415 642494 448455 642814
rect 448055 642454 448455 642494
rect 448774 642814 449174 642854
rect 448774 642494 448814 642814
rect 449134 642494 449174 642814
rect 448774 642454 449174 642494
rect 449493 642814 449893 642854
rect 449493 642494 449533 642814
rect 449853 642494 449893 642814
rect 449493 642454 449893 642494
rect 450212 642814 450612 642854
rect 450212 642494 450252 642814
rect 450572 642494 450612 642814
rect 450212 642454 450612 642494
rect 450931 642814 451331 642854
rect 450931 642494 450971 642814
rect 451291 642494 451331 642814
rect 450931 642454 451331 642494
rect 444460 642114 444860 642154
rect 444460 641794 444500 642114
rect 444820 641794 444860 642114
rect 444460 641754 444860 641794
rect 445179 642114 445579 642154
rect 445179 641794 445219 642114
rect 445539 641794 445579 642114
rect 445179 641754 445579 641794
rect 445898 642114 446298 642154
rect 445898 641794 445938 642114
rect 446258 641794 446298 642114
rect 445898 641754 446298 641794
rect 446617 642114 447017 642154
rect 446617 641794 446657 642114
rect 446977 641794 447017 642114
rect 446617 641754 447017 641794
rect 447336 642114 447736 642154
rect 447336 641794 447376 642114
rect 447696 641794 447736 642114
rect 447336 641754 447736 641794
rect 448055 642114 448455 642154
rect 448055 641794 448095 642114
rect 448415 641794 448455 642114
rect 448055 641754 448455 641794
rect 448774 642114 449174 642154
rect 448774 641794 448814 642114
rect 449134 641794 449174 642114
rect 448774 641754 449174 641794
rect 449493 642114 449893 642154
rect 449493 641794 449533 642114
rect 449853 641794 449893 642114
rect 449493 641754 449893 641794
rect 450212 642114 450612 642154
rect 450212 641794 450252 642114
rect 450572 641794 450612 642114
rect 450212 641754 450612 641794
rect 450931 642114 451331 642154
rect 450931 641794 450971 642114
rect 451291 641794 451331 642114
rect 450931 641754 451331 641794
rect 444460 641414 444860 641454
rect 444460 641094 444500 641414
rect 444820 641094 444860 641414
rect 444460 641054 444860 641094
rect 445179 641414 445579 641454
rect 445179 641094 445219 641414
rect 445539 641094 445579 641414
rect 445179 641054 445579 641094
rect 445898 641414 446298 641454
rect 445898 641094 445938 641414
rect 446258 641094 446298 641414
rect 445898 641054 446298 641094
rect 446617 641414 447017 641454
rect 446617 641094 446657 641414
rect 446977 641094 447017 641414
rect 446617 641054 447017 641094
rect 447336 641414 447736 641454
rect 447336 641094 447376 641414
rect 447696 641094 447736 641414
rect 447336 641054 447736 641094
rect 448055 641414 448455 641454
rect 448055 641094 448095 641414
rect 448415 641094 448455 641414
rect 448055 641054 448455 641094
rect 448774 641414 449174 641454
rect 448774 641094 448814 641414
rect 449134 641094 449174 641414
rect 448774 641054 449174 641094
rect 449493 641414 449893 641454
rect 449493 641094 449533 641414
rect 449853 641094 449893 641414
rect 449493 641054 449893 641094
rect 450212 641414 450612 641454
rect 450212 641094 450252 641414
rect 450572 641094 450612 641414
rect 450212 641054 450612 641094
rect 450931 641414 451331 641454
rect 450931 641094 450971 641414
rect 451291 641094 451331 641414
rect 450931 641054 451331 641094
rect 444460 640714 444860 640754
rect 444460 640394 444500 640714
rect 444820 640394 444860 640714
rect 444460 640354 444860 640394
rect 445179 640714 445579 640754
rect 445179 640394 445219 640714
rect 445539 640394 445579 640714
rect 445179 640354 445579 640394
rect 445898 640714 446298 640754
rect 445898 640394 445938 640714
rect 446258 640394 446298 640714
rect 445898 640354 446298 640394
rect 446617 640714 447017 640754
rect 446617 640394 446657 640714
rect 446977 640394 447017 640714
rect 446617 640354 447017 640394
rect 447336 640714 447736 640754
rect 447336 640394 447376 640714
rect 447696 640394 447736 640714
rect 447336 640354 447736 640394
rect 448055 640714 448455 640754
rect 448055 640394 448095 640714
rect 448415 640394 448455 640714
rect 448055 640354 448455 640394
rect 448774 640714 449174 640754
rect 448774 640394 448814 640714
rect 449134 640394 449174 640714
rect 448774 640354 449174 640394
rect 449493 640714 449893 640754
rect 449493 640394 449533 640714
rect 449853 640394 449893 640714
rect 449493 640354 449893 640394
rect 450212 640714 450612 640754
rect 450212 640394 450252 640714
rect 450572 640394 450612 640714
rect 450212 640354 450612 640394
rect 450931 640714 451331 640754
rect 450931 640394 450971 640714
rect 451291 640394 451331 640714
rect 450931 640354 451331 640394
rect 444460 640014 444860 640054
rect 444460 639694 444500 640014
rect 444820 639694 444860 640014
rect 444460 639654 444860 639694
rect 445179 640014 445579 640054
rect 445179 639694 445219 640014
rect 445539 639694 445579 640014
rect 445179 639654 445579 639694
rect 445898 640014 446298 640054
rect 445898 639694 445938 640014
rect 446258 639694 446298 640014
rect 445898 639654 446298 639694
rect 446617 640014 447017 640054
rect 446617 639694 446657 640014
rect 446977 639694 447017 640014
rect 446617 639654 447017 639694
rect 447336 640014 447736 640054
rect 447336 639694 447376 640014
rect 447696 639694 447736 640014
rect 447336 639654 447736 639694
rect 448055 640014 448455 640054
rect 448055 639694 448095 640014
rect 448415 639694 448455 640014
rect 448055 639654 448455 639694
rect 448774 640014 449174 640054
rect 448774 639694 448814 640014
rect 449134 639694 449174 640014
rect 448774 639654 449174 639694
rect 449493 640014 449893 640054
rect 449493 639694 449533 640014
rect 449853 639694 449893 640014
rect 449493 639654 449893 639694
rect 450212 640014 450612 640054
rect 450212 639694 450252 640014
rect 450572 639694 450612 640014
rect 450212 639654 450612 639694
rect 450931 640014 451331 640054
rect 450931 639694 450971 640014
rect 451291 639694 451331 640014
rect 450931 639654 451331 639694
rect 444460 639314 444860 639354
rect 444460 638994 444500 639314
rect 444820 638994 444860 639314
rect 444460 638954 444860 638994
rect 445179 639314 445579 639354
rect 445179 638994 445219 639314
rect 445539 638994 445579 639314
rect 445179 638954 445579 638994
rect 445898 639314 446298 639354
rect 445898 638994 445938 639314
rect 446258 638994 446298 639314
rect 445898 638954 446298 638994
rect 446617 639314 447017 639354
rect 446617 638994 446657 639314
rect 446977 638994 447017 639314
rect 446617 638954 447017 638994
rect 447336 639314 447736 639354
rect 447336 638994 447376 639314
rect 447696 638994 447736 639314
rect 447336 638954 447736 638994
rect 448055 639314 448455 639354
rect 448055 638994 448095 639314
rect 448415 638994 448455 639314
rect 448055 638954 448455 638994
rect 448774 639314 449174 639354
rect 448774 638994 448814 639314
rect 449134 638994 449174 639314
rect 448774 638954 449174 638994
rect 449493 639314 449893 639354
rect 449493 638994 449533 639314
rect 449853 638994 449893 639314
rect 449493 638954 449893 638994
rect 450212 639314 450612 639354
rect 450212 638994 450252 639314
rect 450572 638994 450612 639314
rect 450212 638954 450612 638994
rect 450931 639314 451331 639354
rect 450931 638994 450971 639314
rect 451291 638994 451331 639314
rect 450931 638954 451331 638994
rect 444460 638614 444860 638654
rect 444460 638294 444500 638614
rect 444820 638294 444860 638614
rect 444460 638254 444860 638294
rect 445179 638614 445579 638654
rect 445179 638294 445219 638614
rect 445539 638294 445579 638614
rect 445179 638254 445579 638294
rect 445898 638614 446298 638654
rect 445898 638294 445938 638614
rect 446258 638294 446298 638614
rect 445898 638254 446298 638294
rect 446617 638614 447017 638654
rect 446617 638294 446657 638614
rect 446977 638294 447017 638614
rect 446617 638254 447017 638294
rect 447336 638614 447736 638654
rect 447336 638294 447376 638614
rect 447696 638294 447736 638614
rect 447336 638254 447736 638294
rect 448055 638614 448455 638654
rect 448055 638294 448095 638614
rect 448415 638294 448455 638614
rect 448055 638254 448455 638294
rect 448774 638614 449174 638654
rect 448774 638294 448814 638614
rect 449134 638294 449174 638614
rect 448774 638254 449174 638294
rect 449493 638614 449893 638654
rect 449493 638294 449533 638614
rect 449853 638294 449893 638614
rect 449493 638254 449893 638294
rect 450212 638614 450612 638654
rect 450212 638294 450252 638614
rect 450572 638294 450612 638614
rect 450212 638254 450612 638294
rect 450931 638614 451331 638654
rect 450931 638294 450971 638614
rect 451291 638294 451331 638614
rect 450931 638254 451331 638294
rect 444460 637914 444860 637954
rect 444460 637594 444500 637914
rect 444820 637594 444860 637914
rect 444460 637554 444860 637594
rect 445179 637914 445579 637954
rect 445179 637594 445219 637914
rect 445539 637594 445579 637914
rect 445179 637554 445579 637594
rect 445898 637914 446298 637954
rect 445898 637594 445938 637914
rect 446258 637594 446298 637914
rect 445898 637554 446298 637594
rect 446617 637914 447017 637954
rect 446617 637594 446657 637914
rect 446977 637594 447017 637914
rect 446617 637554 447017 637594
rect 447336 637914 447736 637954
rect 447336 637594 447376 637914
rect 447696 637594 447736 637914
rect 447336 637554 447736 637594
rect 448055 637914 448455 637954
rect 448055 637594 448095 637914
rect 448415 637594 448455 637914
rect 448055 637554 448455 637594
rect 448774 637914 449174 637954
rect 448774 637594 448814 637914
rect 449134 637594 449174 637914
rect 448774 637554 449174 637594
rect 449493 637914 449893 637954
rect 449493 637594 449533 637914
rect 449853 637594 449893 637914
rect 449493 637554 449893 637594
rect 450212 637914 450612 637954
rect 450212 637594 450252 637914
rect 450572 637594 450612 637914
rect 450212 637554 450612 637594
rect 450931 637914 451331 637954
rect 450931 637594 450971 637914
rect 451291 637594 451331 637914
rect 450931 637554 451331 637594
<< mimcapcontact >>
rect 444500 643894 444820 644214
rect 445219 643894 445539 644214
rect 445938 643894 446258 644214
rect 446657 643894 446977 644214
rect 447376 643894 447696 644214
rect 448095 643894 448415 644214
rect 448814 643894 449134 644214
rect 449533 643894 449853 644214
rect 450252 643894 450572 644214
rect 450971 643894 451291 644214
rect 444500 643194 444820 643514
rect 445219 643194 445539 643514
rect 445938 643194 446258 643514
rect 446657 643194 446977 643514
rect 447376 643194 447696 643514
rect 448095 643194 448415 643514
rect 448814 643194 449134 643514
rect 449533 643194 449853 643514
rect 450252 643194 450572 643514
rect 450971 643194 451291 643514
rect 444500 642494 444820 642814
rect 445219 642494 445539 642814
rect 445938 642494 446258 642814
rect 446657 642494 446977 642814
rect 447376 642494 447696 642814
rect 448095 642494 448415 642814
rect 448814 642494 449134 642814
rect 449533 642494 449853 642814
rect 450252 642494 450572 642814
rect 450971 642494 451291 642814
rect 444500 641794 444820 642114
rect 445219 641794 445539 642114
rect 445938 641794 446258 642114
rect 446657 641794 446977 642114
rect 447376 641794 447696 642114
rect 448095 641794 448415 642114
rect 448814 641794 449134 642114
rect 449533 641794 449853 642114
rect 450252 641794 450572 642114
rect 450971 641794 451291 642114
rect 444500 641094 444820 641414
rect 445219 641094 445539 641414
rect 445938 641094 446258 641414
rect 446657 641094 446977 641414
rect 447376 641094 447696 641414
rect 448095 641094 448415 641414
rect 448814 641094 449134 641414
rect 449533 641094 449853 641414
rect 450252 641094 450572 641414
rect 450971 641094 451291 641414
rect 444500 640394 444820 640714
rect 445219 640394 445539 640714
rect 445938 640394 446258 640714
rect 446657 640394 446977 640714
rect 447376 640394 447696 640714
rect 448095 640394 448415 640714
rect 448814 640394 449134 640714
rect 449533 640394 449853 640714
rect 450252 640394 450572 640714
rect 450971 640394 451291 640714
rect 444500 639694 444820 640014
rect 445219 639694 445539 640014
rect 445938 639694 446258 640014
rect 446657 639694 446977 640014
rect 447376 639694 447696 640014
rect 448095 639694 448415 640014
rect 448814 639694 449134 640014
rect 449533 639694 449853 640014
rect 450252 639694 450572 640014
rect 450971 639694 451291 640014
rect 444500 638994 444820 639314
rect 445219 638994 445539 639314
rect 445938 638994 446258 639314
rect 446657 638994 446977 639314
rect 447376 638994 447696 639314
rect 448095 638994 448415 639314
rect 448814 638994 449134 639314
rect 449533 638994 449853 639314
rect 450252 638994 450572 639314
rect 450971 638994 451291 639314
rect 444500 638294 444820 638614
rect 445219 638294 445539 638614
rect 445938 638294 446258 638614
rect 446657 638294 446977 638614
rect 447376 638294 447696 638614
rect 448095 638294 448415 638614
rect 448814 638294 449134 638614
rect 449533 638294 449853 638614
rect 450252 638294 450572 638614
rect 450971 638294 451291 638614
rect 444500 637594 444820 637914
rect 445219 637594 445539 637914
rect 445938 637594 446258 637914
rect 446657 637594 446977 637914
rect 447376 637594 447696 637914
rect 448095 637594 448415 637914
rect 448814 637594 449134 637914
rect 449533 637594 449853 637914
rect 450252 637594 450572 637914
rect 450971 637594 451291 637914
<< metal4 >>
rect 483464 663582 487922 663588
rect 425844 663144 497922 663582
rect 425844 663086 487200 663144
rect 425844 662766 476524 663086
rect 425844 657022 429964 662766
rect 434748 657022 438964 662766
rect 443748 657022 444964 662766
rect 449748 657022 450964 662766
rect 455748 657342 476524 662766
rect 481308 657400 487200 663086
rect 491984 657400 497922 663144
rect 481308 657342 497922 657400
rect 455748 657022 497922 657342
rect 425844 656926 497922 657022
rect 475604 654901 482260 654906
rect 475604 654896 482261 654901
rect 438864 654881 445520 654886
rect 449334 654881 455990 654886
rect 438864 654876 445521 654881
rect 438864 654776 438920 654876
rect 439020 654776 439144 654876
rect 439244 654776 439368 654876
rect 439468 654776 439592 654876
rect 439692 654776 439816 654876
rect 439916 654776 440040 654876
rect 440140 654776 440264 654876
rect 440364 654776 440488 654876
rect 440588 654776 440712 654876
rect 440812 654776 440936 654876
rect 441036 654776 441160 654876
rect 441260 654776 441384 654876
rect 441484 654776 441608 654876
rect 441708 654776 441832 654876
rect 441932 654776 442056 654876
rect 442156 654776 442280 654876
rect 442380 654776 442504 654876
rect 442604 654776 442728 654876
rect 442828 654776 442952 654876
rect 443052 654776 443176 654876
rect 443276 654776 443400 654876
rect 443500 654776 443624 654876
rect 443724 654776 443848 654876
rect 443948 654776 444072 654876
rect 444172 654776 444296 654876
rect 444396 654776 444520 654876
rect 444620 654776 444744 654876
rect 444844 654776 444968 654876
rect 445068 654776 445192 654876
rect 445292 654776 445416 654876
rect 445516 654776 445521 654876
rect 438864 654771 445521 654776
rect 449334 654876 455991 654881
rect 449334 654776 449390 654876
rect 449490 654776 449614 654876
rect 449714 654776 449838 654876
rect 449938 654776 450062 654876
rect 450162 654776 450286 654876
rect 450386 654776 450510 654876
rect 450610 654776 450734 654876
rect 450834 654776 450958 654876
rect 451058 654776 451182 654876
rect 451282 654776 451406 654876
rect 451506 654776 451630 654876
rect 451730 654776 451854 654876
rect 451954 654776 452078 654876
rect 452178 654776 452302 654876
rect 452402 654776 452526 654876
rect 452626 654776 452750 654876
rect 452850 654776 452974 654876
rect 453074 654776 453198 654876
rect 453298 654776 453422 654876
rect 453522 654776 453646 654876
rect 453746 654776 453870 654876
rect 453970 654776 454094 654876
rect 454194 654776 454318 654876
rect 454418 654776 454542 654876
rect 454642 654776 454766 654876
rect 454866 654776 454990 654876
rect 455090 654776 455214 654876
rect 455314 654776 455438 654876
rect 455538 654776 455662 654876
rect 455762 654776 455886 654876
rect 455986 654776 455991 654876
rect 449334 654771 455991 654776
rect 475604 654796 475660 654896
rect 475760 654796 475884 654896
rect 475984 654796 476108 654896
rect 476208 654796 476332 654896
rect 476432 654796 476556 654896
rect 476656 654796 476780 654896
rect 476880 654796 477004 654896
rect 477104 654796 477228 654896
rect 477328 654796 477452 654896
rect 477552 654796 477676 654896
rect 477776 654796 477900 654896
rect 478000 654796 478124 654896
rect 478224 654796 478348 654896
rect 478448 654796 478572 654896
rect 478672 654796 478796 654896
rect 478896 654796 479020 654896
rect 479120 654796 479244 654896
rect 479344 654796 479468 654896
rect 479568 654796 479692 654896
rect 479792 654796 479916 654896
rect 480016 654796 480140 654896
rect 480240 654796 480364 654896
rect 480464 654796 480588 654896
rect 480688 654796 480812 654896
rect 480912 654796 481036 654896
rect 481136 654796 481260 654896
rect 481360 654796 481484 654896
rect 481584 654796 481708 654896
rect 481808 654796 481932 654896
rect 482032 654796 482156 654896
rect 482256 654796 482261 654896
rect 475604 654791 482261 654796
rect 438864 654657 445520 654771
rect 449334 654657 455990 654771
rect 475604 654677 482260 654791
rect 475604 654672 482261 654677
rect 438864 654652 445521 654657
rect 438864 654552 438920 654652
rect 439020 654552 439144 654652
rect 439244 654552 439368 654652
rect 439468 654552 439592 654652
rect 439692 654552 439816 654652
rect 439916 654552 440040 654652
rect 440140 654552 440264 654652
rect 440364 654552 440488 654652
rect 440588 654552 440712 654652
rect 440812 654552 440936 654652
rect 441036 654552 441160 654652
rect 441260 654552 441384 654652
rect 441484 654552 441608 654652
rect 441708 654552 441832 654652
rect 441932 654552 442056 654652
rect 442156 654552 442280 654652
rect 442380 654552 442504 654652
rect 442604 654552 442728 654652
rect 442828 654552 442952 654652
rect 443052 654552 443176 654652
rect 443276 654552 443400 654652
rect 443500 654552 443624 654652
rect 443724 654552 443848 654652
rect 443948 654552 444072 654652
rect 444172 654552 444296 654652
rect 444396 654552 444520 654652
rect 444620 654552 444744 654652
rect 444844 654552 444968 654652
rect 445068 654552 445192 654652
rect 445292 654552 445416 654652
rect 445516 654552 445521 654652
rect 438864 654547 445521 654552
rect 449334 654652 455991 654657
rect 449334 654552 449390 654652
rect 449490 654552 449614 654652
rect 449714 654552 449838 654652
rect 449938 654552 450062 654652
rect 450162 654552 450286 654652
rect 450386 654552 450510 654652
rect 450610 654552 450734 654652
rect 450834 654552 450958 654652
rect 451058 654552 451182 654652
rect 451282 654552 451406 654652
rect 451506 654552 451630 654652
rect 451730 654552 451854 654652
rect 451954 654552 452078 654652
rect 452178 654552 452302 654652
rect 452402 654552 452526 654652
rect 452626 654552 452750 654652
rect 452850 654552 452974 654652
rect 453074 654552 453198 654652
rect 453298 654552 453422 654652
rect 453522 654552 453646 654652
rect 453746 654552 453870 654652
rect 453970 654552 454094 654652
rect 454194 654552 454318 654652
rect 454418 654552 454542 654652
rect 454642 654552 454766 654652
rect 454866 654552 454990 654652
rect 455090 654552 455214 654652
rect 455314 654552 455438 654652
rect 455538 654552 455662 654652
rect 455762 654552 455886 654652
rect 455986 654552 455991 654652
rect 449334 654547 455991 654552
rect 475604 654572 475660 654672
rect 475760 654572 475884 654672
rect 475984 654572 476108 654672
rect 476208 654572 476332 654672
rect 476432 654572 476556 654672
rect 476656 654572 476780 654672
rect 476880 654572 477004 654672
rect 477104 654572 477228 654672
rect 477328 654572 477452 654672
rect 477552 654572 477676 654672
rect 477776 654572 477900 654672
rect 478000 654572 478124 654672
rect 478224 654572 478348 654672
rect 478448 654572 478572 654672
rect 478672 654572 478796 654672
rect 478896 654572 479020 654672
rect 479120 654572 479244 654672
rect 479344 654572 479468 654672
rect 479568 654572 479692 654672
rect 479792 654572 479916 654672
rect 480016 654572 480140 654672
rect 480240 654572 480364 654672
rect 480464 654572 480588 654672
rect 480688 654572 480812 654672
rect 480912 654572 481036 654672
rect 481136 654572 481260 654672
rect 481360 654572 481484 654672
rect 481584 654572 481708 654672
rect 481808 654572 481932 654672
rect 482032 654572 482156 654672
rect 482256 654572 482261 654672
rect 475604 654567 482261 654572
rect 438864 654433 445520 654547
rect 449334 654433 455990 654547
rect 475604 654453 482260 654567
rect 475604 654448 482261 654453
rect 438864 654428 445521 654433
rect 438864 654328 438920 654428
rect 439020 654328 439144 654428
rect 439244 654328 439368 654428
rect 439468 654328 439592 654428
rect 439692 654328 439816 654428
rect 439916 654328 440040 654428
rect 440140 654328 440264 654428
rect 440364 654328 440488 654428
rect 440588 654328 440712 654428
rect 440812 654328 440936 654428
rect 441036 654328 441160 654428
rect 441260 654328 441384 654428
rect 441484 654328 441608 654428
rect 441708 654328 441832 654428
rect 441932 654328 442056 654428
rect 442156 654328 442280 654428
rect 442380 654328 442504 654428
rect 442604 654328 442728 654428
rect 442828 654328 442952 654428
rect 443052 654328 443176 654428
rect 443276 654328 443400 654428
rect 443500 654328 443624 654428
rect 443724 654328 443848 654428
rect 443948 654328 444072 654428
rect 444172 654328 444296 654428
rect 444396 654328 444520 654428
rect 444620 654328 444744 654428
rect 444844 654328 444968 654428
rect 445068 654328 445192 654428
rect 445292 654328 445416 654428
rect 445516 654328 445521 654428
rect 438864 654323 445521 654328
rect 449334 654428 455991 654433
rect 449334 654328 449390 654428
rect 449490 654328 449614 654428
rect 449714 654328 449838 654428
rect 449938 654328 450062 654428
rect 450162 654328 450286 654428
rect 450386 654328 450510 654428
rect 450610 654328 450734 654428
rect 450834 654328 450958 654428
rect 451058 654328 451182 654428
rect 451282 654328 451406 654428
rect 451506 654328 451630 654428
rect 451730 654328 451854 654428
rect 451954 654328 452078 654428
rect 452178 654328 452302 654428
rect 452402 654328 452526 654428
rect 452626 654328 452750 654428
rect 452850 654328 452974 654428
rect 453074 654328 453198 654428
rect 453298 654328 453422 654428
rect 453522 654328 453646 654428
rect 453746 654328 453870 654428
rect 453970 654328 454094 654428
rect 454194 654328 454318 654428
rect 454418 654328 454542 654428
rect 454642 654328 454766 654428
rect 454866 654328 454990 654428
rect 455090 654328 455214 654428
rect 455314 654328 455438 654428
rect 455538 654328 455662 654428
rect 455762 654328 455886 654428
rect 455986 654328 455991 654428
rect 449334 654323 455991 654328
rect 475604 654348 475660 654448
rect 475760 654348 475884 654448
rect 475984 654348 476108 654448
rect 476208 654348 476332 654448
rect 476432 654348 476556 654448
rect 476656 654348 476780 654448
rect 476880 654348 477004 654448
rect 477104 654348 477228 654448
rect 477328 654348 477452 654448
rect 477552 654348 477676 654448
rect 477776 654348 477900 654448
rect 478000 654348 478124 654448
rect 478224 654348 478348 654448
rect 478448 654348 478572 654448
rect 478672 654348 478796 654448
rect 478896 654348 479020 654448
rect 479120 654348 479244 654448
rect 479344 654348 479468 654448
rect 479568 654348 479692 654448
rect 479792 654348 479916 654448
rect 480016 654348 480140 654448
rect 480240 654348 480364 654448
rect 480464 654348 480588 654448
rect 480688 654348 480812 654448
rect 480912 654348 481036 654448
rect 481136 654348 481260 654448
rect 481360 654348 481484 654448
rect 481584 654348 481708 654448
rect 481808 654348 481932 654448
rect 482032 654348 482156 654448
rect 482256 654348 482261 654448
rect 475604 654343 482261 654348
rect 438864 654209 445520 654323
rect 449334 654209 455990 654323
rect 475604 654229 482260 654343
rect 475604 654224 482261 654229
rect 438864 654204 445521 654209
rect 438864 654104 438920 654204
rect 439020 654104 439144 654204
rect 439244 654104 439368 654204
rect 439468 654104 439592 654204
rect 439692 654104 439816 654204
rect 439916 654104 440040 654204
rect 440140 654104 440264 654204
rect 440364 654104 440488 654204
rect 440588 654104 440712 654204
rect 440812 654104 440936 654204
rect 441036 654104 441160 654204
rect 441260 654104 441384 654204
rect 441484 654104 441608 654204
rect 441708 654104 441832 654204
rect 441932 654104 442056 654204
rect 442156 654104 442280 654204
rect 442380 654104 442504 654204
rect 442604 654104 442728 654204
rect 442828 654104 442952 654204
rect 443052 654104 443176 654204
rect 443276 654104 443400 654204
rect 443500 654104 443624 654204
rect 443724 654104 443848 654204
rect 443948 654104 444072 654204
rect 444172 654104 444296 654204
rect 444396 654104 444520 654204
rect 444620 654104 444744 654204
rect 444844 654104 444968 654204
rect 445068 654104 445192 654204
rect 445292 654104 445416 654204
rect 445516 654104 445521 654204
rect 438864 654099 445521 654104
rect 449334 654204 455991 654209
rect 449334 654104 449390 654204
rect 449490 654104 449614 654204
rect 449714 654104 449838 654204
rect 449938 654104 450062 654204
rect 450162 654104 450286 654204
rect 450386 654104 450510 654204
rect 450610 654104 450734 654204
rect 450834 654104 450958 654204
rect 451058 654104 451182 654204
rect 451282 654104 451406 654204
rect 451506 654104 451630 654204
rect 451730 654104 451854 654204
rect 451954 654104 452078 654204
rect 452178 654104 452302 654204
rect 452402 654104 452526 654204
rect 452626 654104 452750 654204
rect 452850 654104 452974 654204
rect 453074 654104 453198 654204
rect 453298 654104 453422 654204
rect 453522 654104 453646 654204
rect 453746 654104 453870 654204
rect 453970 654104 454094 654204
rect 454194 654104 454318 654204
rect 454418 654104 454542 654204
rect 454642 654104 454766 654204
rect 454866 654104 454990 654204
rect 455090 654104 455214 654204
rect 455314 654104 455438 654204
rect 455538 654104 455662 654204
rect 455762 654104 455886 654204
rect 455986 654104 455991 654204
rect 449334 654099 455991 654104
rect 475604 654124 475660 654224
rect 475760 654124 475884 654224
rect 475984 654124 476108 654224
rect 476208 654124 476332 654224
rect 476432 654124 476556 654224
rect 476656 654124 476780 654224
rect 476880 654124 477004 654224
rect 477104 654124 477228 654224
rect 477328 654124 477452 654224
rect 477552 654124 477676 654224
rect 477776 654124 477900 654224
rect 478000 654124 478124 654224
rect 478224 654124 478348 654224
rect 478448 654124 478572 654224
rect 478672 654124 478796 654224
rect 478896 654124 479020 654224
rect 479120 654124 479244 654224
rect 479344 654124 479468 654224
rect 479568 654124 479692 654224
rect 479792 654124 479916 654224
rect 480016 654124 480140 654224
rect 480240 654124 480364 654224
rect 480464 654124 480588 654224
rect 480688 654124 480812 654224
rect 480912 654124 481036 654224
rect 481136 654124 481260 654224
rect 481360 654124 481484 654224
rect 481584 654124 481708 654224
rect 481808 654124 481932 654224
rect 482032 654124 482156 654224
rect 482256 654124 482261 654224
rect 475604 654119 482261 654124
rect 438864 653985 445520 654099
rect 449334 653985 455990 654099
rect 475604 654005 482260 654119
rect 475604 654000 482261 654005
rect 438864 653980 445521 653985
rect 438864 653880 438920 653980
rect 439020 653880 439144 653980
rect 439244 653880 439368 653980
rect 439468 653880 439592 653980
rect 439692 653880 439816 653980
rect 439916 653880 440040 653980
rect 440140 653880 440264 653980
rect 440364 653880 440488 653980
rect 440588 653880 440712 653980
rect 440812 653880 440936 653980
rect 441036 653880 441160 653980
rect 441260 653880 441384 653980
rect 441484 653880 441608 653980
rect 441708 653880 441832 653980
rect 441932 653880 442056 653980
rect 442156 653880 442280 653980
rect 442380 653880 442504 653980
rect 442604 653880 442728 653980
rect 442828 653880 442952 653980
rect 443052 653880 443176 653980
rect 443276 653880 443400 653980
rect 443500 653880 443624 653980
rect 443724 653880 443848 653980
rect 443948 653880 444072 653980
rect 444172 653880 444296 653980
rect 444396 653880 444520 653980
rect 444620 653880 444744 653980
rect 444844 653880 444968 653980
rect 445068 653880 445192 653980
rect 445292 653880 445416 653980
rect 445516 653880 445521 653980
rect 438864 653875 445521 653880
rect 449334 653980 455991 653985
rect 449334 653880 449390 653980
rect 449490 653880 449614 653980
rect 449714 653880 449838 653980
rect 449938 653880 450062 653980
rect 450162 653880 450286 653980
rect 450386 653880 450510 653980
rect 450610 653880 450734 653980
rect 450834 653880 450958 653980
rect 451058 653880 451182 653980
rect 451282 653880 451406 653980
rect 451506 653880 451630 653980
rect 451730 653880 451854 653980
rect 451954 653880 452078 653980
rect 452178 653880 452302 653980
rect 452402 653880 452526 653980
rect 452626 653880 452750 653980
rect 452850 653880 452974 653980
rect 453074 653880 453198 653980
rect 453298 653880 453422 653980
rect 453522 653880 453646 653980
rect 453746 653880 453870 653980
rect 453970 653880 454094 653980
rect 454194 653880 454318 653980
rect 454418 653880 454542 653980
rect 454642 653880 454766 653980
rect 454866 653880 454990 653980
rect 455090 653880 455214 653980
rect 455314 653880 455438 653980
rect 455538 653880 455662 653980
rect 455762 653880 455886 653980
rect 455986 653880 455991 653980
rect 449334 653875 455991 653880
rect 475604 653900 475660 654000
rect 475760 653900 475884 654000
rect 475984 653900 476108 654000
rect 476208 653900 476332 654000
rect 476432 653900 476556 654000
rect 476656 653900 476780 654000
rect 476880 653900 477004 654000
rect 477104 653900 477228 654000
rect 477328 653900 477452 654000
rect 477552 653900 477676 654000
rect 477776 653900 477900 654000
rect 478000 653900 478124 654000
rect 478224 653900 478348 654000
rect 478448 653900 478572 654000
rect 478672 653900 478796 654000
rect 478896 653900 479020 654000
rect 479120 653900 479244 654000
rect 479344 653900 479468 654000
rect 479568 653900 479692 654000
rect 479792 653900 479916 654000
rect 480016 653900 480140 654000
rect 480240 653900 480364 654000
rect 480464 653900 480588 654000
rect 480688 653900 480812 654000
rect 480912 653900 481036 654000
rect 481136 653900 481260 654000
rect 481360 653900 481484 654000
rect 481584 653900 481708 654000
rect 481808 653900 481932 654000
rect 482032 653900 482156 654000
rect 482256 653900 482261 654000
rect 475604 653895 482261 653900
rect 438864 653846 445520 653875
rect 449334 653846 455990 653875
rect 475604 653866 482260 653895
rect 440670 652769 451996 652806
rect 440670 651913 440687 652769
rect 451961 651913 451996 652769
rect 429064 650178 438924 650202
rect 429064 650078 437894 650178
rect 437994 650078 438118 650178
rect 438218 650078 438342 650178
rect 438442 650078 438566 650178
rect 438666 650078 438790 650178
rect 438890 650078 438924 650178
rect 429064 649954 438924 650078
rect 429064 649854 437894 649954
rect 437994 649854 438118 649954
rect 438218 649854 438342 649954
rect 438442 649854 438566 649954
rect 438666 649854 438790 649954
rect 438890 649854 438924 649954
rect 429064 649730 438924 649854
rect 429064 649630 437894 649730
rect 437994 649630 438118 649730
rect 438218 649630 438342 649730
rect 438442 649630 438566 649730
rect 438666 649630 438790 649730
rect 438890 649630 438924 649730
rect 429064 649506 438924 649630
rect 429064 649406 437894 649506
rect 437994 649406 438118 649506
rect 438218 649406 438342 649506
rect 438442 649406 438566 649506
rect 438666 649406 438790 649506
rect 438890 649406 438924 649506
rect 429064 649366 438924 649406
rect 429064 643622 429964 649366
rect 434748 649282 438924 649366
rect 434748 649182 437894 649282
rect 437994 649182 438118 649282
rect 438218 649182 438342 649282
rect 438442 649182 438566 649282
rect 438666 649182 438790 649282
rect 438890 649182 438924 649282
rect 434748 649058 438924 649182
rect 434748 648958 437894 649058
rect 437994 648958 438118 649058
rect 438218 648958 438342 649058
rect 438442 648958 438566 649058
rect 438666 648958 438790 649058
rect 438890 648958 438924 649058
rect 434748 648834 438924 648958
rect 434748 648734 437894 648834
rect 437994 648734 438118 648834
rect 438218 648734 438342 648834
rect 438442 648734 438566 648834
rect 438666 648734 438790 648834
rect 438890 648734 438924 648834
rect 434748 648610 438924 648734
rect 434748 648510 437894 648610
rect 437994 648510 438118 648610
rect 438218 648510 438342 648610
rect 438442 648510 438566 648610
rect 438666 648510 438790 648610
rect 438890 648510 438924 648610
rect 434748 648386 438924 648510
rect 434748 648286 437894 648386
rect 437994 648286 438118 648386
rect 438218 648286 438342 648386
rect 438442 648286 438566 648386
rect 438666 648286 438790 648386
rect 438890 648286 438924 648386
rect 434748 648162 438924 648286
rect 434748 648062 437894 648162
rect 437994 648062 438118 648162
rect 438218 648062 438342 648162
rect 438442 648062 438566 648162
rect 438666 648062 438790 648162
rect 438890 648062 438924 648162
rect 434748 647938 438924 648062
rect 434748 647838 437894 647938
rect 437994 647838 438118 647938
rect 438218 647838 438342 647938
rect 438442 647838 438566 647938
rect 438666 647838 438790 647938
rect 438890 647838 438924 647938
rect 434748 647714 438924 647838
rect 434748 647614 437894 647714
rect 437994 647614 438118 647714
rect 438218 647614 438342 647714
rect 438442 647614 438566 647714
rect 438666 647614 438790 647714
rect 438890 647614 438924 647714
rect 434748 647490 438924 647614
rect 434748 647390 437894 647490
rect 437994 647390 438118 647490
rect 438218 647390 438342 647490
rect 438442 647390 438566 647490
rect 438666 647390 438790 647490
rect 438890 647390 438924 647490
rect 434748 647266 438924 647390
rect 434748 647166 437894 647266
rect 437994 647166 438118 647266
rect 438218 647166 438342 647266
rect 438442 647166 438566 647266
rect 438666 647166 438790 647266
rect 438890 647166 438924 647266
rect 434748 647042 438924 647166
rect 434748 646942 437894 647042
rect 437994 646942 438118 647042
rect 438218 646942 438342 647042
rect 438442 646942 438566 647042
rect 438666 646942 438790 647042
rect 438890 646942 438924 647042
rect 434748 646818 438924 646942
rect 434748 646718 437894 646818
rect 437994 646718 438118 646818
rect 438218 646718 438342 646818
rect 438442 646718 438566 646818
rect 438666 646718 438790 646818
rect 438890 646718 438924 646818
rect 434748 646594 438924 646718
rect 434748 646494 437894 646594
rect 437994 646494 438118 646594
rect 438218 646494 438342 646594
rect 438442 646494 438566 646594
rect 438666 646494 438790 646594
rect 438890 646494 438924 646594
rect 434748 646370 438924 646494
rect 434748 646270 437894 646370
rect 437994 646270 438118 646370
rect 438218 646270 438342 646370
rect 438442 646270 438566 646370
rect 438666 646270 438790 646370
rect 438890 646270 438924 646370
rect 434748 646146 438924 646270
rect 434748 646046 437894 646146
rect 437994 646046 438118 646146
rect 438218 646046 438342 646146
rect 438442 646046 438566 646146
rect 438666 646046 438790 646146
rect 438890 646046 438924 646146
rect 434748 645922 438924 646046
rect 434748 645822 437894 645922
rect 437994 645822 438118 645922
rect 438218 645822 438342 645922
rect 438442 645822 438566 645922
rect 438666 645822 438790 645922
rect 438890 645822 438924 645922
rect 434748 645698 438924 645822
rect 434748 645598 437894 645698
rect 437994 645598 438118 645698
rect 438218 645598 438342 645698
rect 438442 645598 438566 645698
rect 438666 645598 438790 645698
rect 438890 645598 438924 645698
rect 434748 645474 438924 645598
rect 434748 645374 437894 645474
rect 437994 645374 438118 645474
rect 438218 645374 438342 645474
rect 438442 645374 438566 645474
rect 438666 645374 438790 645474
rect 438890 645374 438924 645474
rect 434748 645250 438924 645374
rect 434748 645150 437894 645250
rect 437994 645150 438118 645250
rect 438218 645150 438342 645250
rect 438442 645150 438566 645250
rect 438666 645150 438790 645250
rect 438890 645150 438924 645250
rect 434748 645026 438924 645150
rect 434748 644926 437894 645026
rect 437994 644926 438118 645026
rect 438218 644926 438342 645026
rect 438442 644926 438566 645026
rect 438666 644926 438790 645026
rect 438890 644926 438924 645026
rect 434748 644802 438924 644926
rect 434748 644702 437894 644802
rect 437994 644702 438118 644802
rect 438218 644702 438342 644802
rect 438442 644702 438566 644802
rect 438666 644702 438790 644802
rect 438890 644702 438924 644802
rect 434748 644578 438924 644702
rect 440670 644644 451996 651913
rect 482169 650182 482279 650183
rect 482393 650182 482503 650183
rect 482617 650182 482727 650183
rect 482841 650182 482951 650183
rect 483065 650182 483175 650183
rect 440716 644638 451996 644644
rect 482038 650178 492674 650182
rect 482038 650078 482174 650178
rect 482274 650078 482398 650178
rect 482498 650078 482622 650178
rect 482722 650078 482846 650178
rect 482946 650078 483070 650178
rect 483170 650078 492674 650178
rect 482038 649954 492674 650078
rect 482038 649854 482174 649954
rect 482274 649854 482398 649954
rect 482498 649854 482622 649954
rect 482722 649854 482846 649954
rect 482946 649854 483070 649954
rect 483170 649854 492674 649954
rect 482038 649744 492674 649854
rect 482038 649730 487200 649744
rect 482038 649630 482174 649730
rect 482274 649630 482398 649730
rect 482498 649630 482622 649730
rect 482722 649630 482846 649730
rect 482946 649630 483070 649730
rect 483170 649630 487200 649730
rect 482038 649506 487200 649630
rect 482038 649406 482174 649506
rect 482274 649406 482398 649506
rect 482498 649406 482622 649506
rect 482722 649406 482846 649506
rect 482946 649406 483070 649506
rect 483170 649406 487200 649506
rect 482038 649282 487200 649406
rect 482038 649182 482174 649282
rect 482274 649182 482398 649282
rect 482498 649182 482622 649282
rect 482722 649182 482846 649282
rect 482946 649182 483070 649282
rect 483170 649182 487200 649282
rect 482038 649058 487200 649182
rect 482038 648958 482174 649058
rect 482274 648958 482398 649058
rect 482498 648958 482622 649058
rect 482722 648958 482846 649058
rect 482946 648958 483070 649058
rect 483170 648958 487200 649058
rect 482038 648834 487200 648958
rect 482038 648734 482174 648834
rect 482274 648734 482398 648834
rect 482498 648734 482622 648834
rect 482722 648734 482846 648834
rect 482946 648734 483070 648834
rect 483170 648734 487200 648834
rect 482038 648610 487200 648734
rect 482038 648510 482174 648610
rect 482274 648510 482398 648610
rect 482498 648510 482622 648610
rect 482722 648510 482846 648610
rect 482946 648510 483070 648610
rect 483170 648510 487200 648610
rect 482038 648386 487200 648510
rect 482038 648286 482174 648386
rect 482274 648286 482398 648386
rect 482498 648286 482622 648386
rect 482722 648286 482846 648386
rect 482946 648286 483070 648386
rect 483170 648286 487200 648386
rect 482038 648162 487200 648286
rect 482038 648062 482174 648162
rect 482274 648062 482398 648162
rect 482498 648062 482622 648162
rect 482722 648062 482846 648162
rect 482946 648062 483070 648162
rect 483170 648062 487200 648162
rect 482038 647938 487200 648062
rect 482038 647838 482174 647938
rect 482274 647838 482398 647938
rect 482498 647838 482622 647938
rect 482722 647838 482846 647938
rect 482946 647838 483070 647938
rect 483170 647838 487200 647938
rect 482038 647714 487200 647838
rect 482038 647614 482174 647714
rect 482274 647614 482398 647714
rect 482498 647614 482622 647714
rect 482722 647614 482846 647714
rect 482946 647614 483070 647714
rect 483170 647614 487200 647714
rect 482038 647490 487200 647614
rect 482038 647390 482174 647490
rect 482274 647390 482398 647490
rect 482498 647390 482622 647490
rect 482722 647390 482846 647490
rect 482946 647390 483070 647490
rect 483170 647390 487200 647490
rect 482038 647266 487200 647390
rect 482038 647166 482174 647266
rect 482274 647166 482398 647266
rect 482498 647166 482622 647266
rect 482722 647166 482846 647266
rect 482946 647166 483070 647266
rect 483170 647166 487200 647266
rect 482038 647042 487200 647166
rect 482038 646942 482174 647042
rect 482274 646942 482398 647042
rect 482498 646942 482622 647042
rect 482722 646942 482846 647042
rect 482946 646942 483070 647042
rect 483170 646942 487200 647042
rect 482038 646818 487200 646942
rect 482038 646718 482174 646818
rect 482274 646718 482398 646818
rect 482498 646718 482622 646818
rect 482722 646718 482846 646818
rect 482946 646718 483070 646818
rect 483170 646718 487200 646818
rect 482038 646594 487200 646718
rect 482038 646494 482174 646594
rect 482274 646494 482398 646594
rect 482498 646494 482622 646594
rect 482722 646494 482846 646594
rect 482946 646494 483070 646594
rect 483170 646494 487200 646594
rect 482038 646370 487200 646494
rect 482038 646270 482174 646370
rect 482274 646270 482398 646370
rect 482498 646270 482622 646370
rect 482722 646270 482846 646370
rect 482946 646270 483070 646370
rect 483170 646270 487200 646370
rect 482038 646146 487200 646270
rect 482038 646046 482174 646146
rect 482274 646046 482398 646146
rect 482498 646046 482622 646146
rect 482722 646046 482846 646146
rect 482946 646046 483070 646146
rect 483170 646046 487200 646146
rect 482038 645922 487200 646046
rect 482038 645822 482174 645922
rect 482274 645822 482398 645922
rect 482498 645822 482622 645922
rect 482722 645822 482846 645922
rect 482946 645822 483070 645922
rect 483170 645822 487200 645922
rect 482038 645698 487200 645822
rect 482038 645598 482174 645698
rect 482274 645598 482398 645698
rect 482498 645598 482622 645698
rect 482722 645598 482846 645698
rect 482946 645598 483070 645698
rect 483170 645598 487200 645698
rect 482038 645474 487200 645598
rect 482038 645374 482174 645474
rect 482274 645374 482398 645474
rect 482498 645374 482622 645474
rect 482722 645374 482846 645474
rect 482946 645374 483070 645474
rect 483170 645374 487200 645474
rect 482038 645250 487200 645374
rect 482038 645150 482174 645250
rect 482274 645150 482398 645250
rect 482498 645150 482622 645250
rect 482722 645150 482846 645250
rect 482946 645150 483070 645250
rect 483170 645150 487200 645250
rect 482038 645026 487200 645150
rect 482038 644926 482174 645026
rect 482274 644926 482398 645026
rect 482498 644926 482622 645026
rect 482722 644926 482846 645026
rect 482946 644926 483070 645026
rect 483170 644926 487200 645026
rect 482038 644802 487200 644926
rect 482038 644702 482174 644802
rect 482274 644702 482398 644802
rect 482498 644702 482622 644802
rect 482722 644702 482846 644802
rect 482946 644702 483070 644802
rect 483170 644702 487200 644802
rect 434748 644478 437894 644578
rect 437994 644478 438118 644578
rect 438218 644478 438342 644578
rect 438442 644478 438566 644578
rect 438666 644478 438790 644578
rect 438890 644478 438924 644578
rect 434748 644354 438924 644478
rect 434748 644254 437894 644354
rect 437994 644254 438118 644354
rect 438218 644254 438342 644354
rect 438442 644254 438566 644354
rect 438666 644254 438790 644354
rect 438890 644254 438924 644354
rect 482038 644578 487200 644702
rect 482038 644478 482174 644578
rect 482274 644478 482398 644578
rect 482498 644478 482622 644578
rect 482722 644478 482846 644578
rect 482946 644478 483070 644578
rect 483170 644478 487200 644578
rect 482038 644354 487200 644478
rect 444959 644326 445055 644342
rect 434748 644130 438924 644254
rect 434748 644030 437894 644130
rect 437994 644030 438118 644130
rect 438218 644030 438342 644130
rect 438442 644030 438566 644130
rect 438666 644030 438790 644130
rect 438890 644030 438924 644130
rect 434748 643906 438924 644030
rect 434748 643806 437894 643906
rect 437994 643806 438118 643906
rect 438218 643806 438342 643906
rect 438442 643806 438566 643906
rect 438666 643806 438790 643906
rect 438890 643806 438924 643906
rect 434748 643682 438924 643806
rect 434748 643622 437894 643682
rect 429064 643582 437894 643622
rect 437994 643582 438118 643682
rect 438218 643582 438342 643682
rect 438442 643582 438566 643682
rect 438666 643582 438790 643682
rect 438890 643582 438924 643682
rect 429064 643522 438924 643582
rect 444460 644214 444860 644254
rect 444460 643894 444500 644214
rect 444820 643894 444860 644214
rect 444460 643514 444860 643894
rect 444959 643782 444975 644326
rect 445039 643782 445055 644326
rect 445678 644326 445774 644342
rect 444959 643766 445055 643782
rect 445180 644214 445580 644254
rect 445180 643894 445219 644214
rect 445539 643894 445580 644214
rect 444460 643194 444500 643514
rect 444820 643194 444860 643514
rect 444460 642814 444860 643194
rect 444959 643626 445055 643642
rect 444959 643082 444975 643626
rect 445039 643082 445055 643626
rect 444959 643066 445055 643082
rect 445180 643514 445580 643894
rect 445678 643782 445694 644326
rect 445758 643782 445774 644326
rect 446397 644326 446493 644342
rect 445678 643766 445774 643782
rect 445900 644214 446300 644254
rect 445900 643894 445938 644214
rect 446258 643894 446300 644214
rect 445180 643194 445219 643514
rect 445539 643194 445580 643514
rect 444460 642494 444500 642814
rect 444820 642494 444860 642814
rect 444460 642114 444860 642494
rect 444959 642926 445055 642942
rect 444959 642382 444975 642926
rect 445039 642382 445055 642926
rect 444959 642366 445055 642382
rect 445180 642814 445580 643194
rect 445678 643626 445774 643642
rect 445678 643082 445694 643626
rect 445758 643082 445774 643626
rect 445678 643066 445774 643082
rect 445900 643514 446300 643894
rect 446397 643782 446413 644326
rect 446477 643782 446493 644326
rect 447116 644326 447212 644342
rect 446397 643766 446493 643782
rect 446620 644214 447020 644254
rect 446620 643894 446657 644214
rect 446977 643894 447020 644214
rect 445900 643194 445938 643514
rect 446258 643194 446300 643514
rect 445180 642494 445219 642814
rect 445539 642494 445580 642814
rect 444460 641794 444500 642114
rect 444820 641794 444860 642114
rect 444460 641414 444860 641794
rect 444959 642226 445055 642242
rect 444959 641682 444975 642226
rect 445039 641682 445055 642226
rect 444959 641666 445055 641682
rect 445180 642114 445580 642494
rect 445678 642926 445774 642942
rect 445678 642382 445694 642926
rect 445758 642382 445774 642926
rect 445678 642366 445774 642382
rect 445900 642814 446300 643194
rect 446397 643626 446493 643642
rect 446397 643082 446413 643626
rect 446477 643082 446493 643626
rect 446397 643066 446493 643082
rect 446620 643514 447020 643894
rect 447116 643782 447132 644326
rect 447196 643782 447212 644326
rect 447835 644326 447931 644342
rect 447116 643766 447212 643782
rect 447340 644214 447740 644254
rect 447340 643894 447376 644214
rect 447696 643894 447740 644214
rect 446620 643194 446657 643514
rect 446977 643194 447020 643514
rect 445900 642494 445938 642814
rect 446258 642494 446300 642814
rect 445180 641794 445219 642114
rect 445539 641794 445580 642114
rect 444460 641094 444500 641414
rect 444820 641094 444860 641414
rect 444460 640714 444860 641094
rect 444959 641526 445055 641542
rect 444959 640982 444975 641526
rect 445039 640982 445055 641526
rect 444959 640966 445055 640982
rect 445180 641414 445580 641794
rect 445678 642226 445774 642242
rect 445678 641682 445694 642226
rect 445758 641682 445774 642226
rect 445678 641666 445774 641682
rect 445900 642114 446300 642494
rect 446397 642926 446493 642942
rect 446397 642382 446413 642926
rect 446477 642382 446493 642926
rect 446397 642366 446493 642382
rect 446620 642814 447020 643194
rect 447116 643626 447212 643642
rect 447116 643082 447132 643626
rect 447196 643082 447212 643626
rect 447116 643066 447212 643082
rect 447340 643514 447740 643894
rect 447835 643782 447851 644326
rect 447915 643782 447931 644326
rect 448554 644326 448650 644342
rect 447835 643766 447931 643782
rect 448060 644214 448460 644254
rect 448060 643894 448095 644214
rect 448415 643894 448460 644214
rect 447340 643194 447376 643514
rect 447696 643194 447740 643514
rect 446620 642494 446657 642814
rect 446977 642494 447020 642814
rect 445900 641794 445938 642114
rect 446258 641794 446300 642114
rect 445180 641094 445219 641414
rect 445539 641094 445580 641414
rect 444460 640394 444500 640714
rect 444820 640394 444860 640714
rect 444460 640014 444860 640394
rect 444959 640826 445055 640842
rect 444959 640282 444975 640826
rect 445039 640282 445055 640826
rect 444959 640266 445055 640282
rect 445180 640714 445580 641094
rect 445678 641526 445774 641542
rect 445678 640982 445694 641526
rect 445758 640982 445774 641526
rect 445678 640966 445774 640982
rect 445900 641414 446300 641794
rect 446397 642226 446493 642242
rect 446397 641682 446413 642226
rect 446477 641682 446493 642226
rect 446397 641666 446493 641682
rect 446620 642114 447020 642494
rect 447116 642926 447212 642942
rect 447116 642382 447132 642926
rect 447196 642382 447212 642926
rect 447116 642366 447212 642382
rect 447340 642814 447740 643194
rect 447835 643626 447931 643642
rect 447835 643082 447851 643626
rect 447915 643082 447931 643626
rect 447835 643066 447931 643082
rect 448060 643514 448460 643894
rect 448554 643782 448570 644326
rect 448634 643782 448650 644326
rect 449273 644326 449369 644342
rect 448554 643766 448650 643782
rect 448780 644214 449180 644254
rect 448780 643894 448814 644214
rect 449134 643894 449180 644214
rect 448060 643194 448095 643514
rect 448415 643194 448460 643514
rect 447340 642494 447376 642814
rect 447696 642494 447740 642814
rect 446620 641794 446657 642114
rect 446977 641794 447020 642114
rect 445900 641094 445938 641414
rect 446258 641094 446300 641414
rect 445180 640394 445219 640714
rect 445539 640394 445580 640714
rect 444460 639694 444500 640014
rect 444820 639694 444860 640014
rect 444460 639314 444860 639694
rect 444959 640126 445055 640142
rect 444959 639582 444975 640126
rect 445039 639582 445055 640126
rect 444959 639566 445055 639582
rect 445180 640014 445580 640394
rect 445678 640826 445774 640842
rect 445678 640282 445694 640826
rect 445758 640282 445774 640826
rect 445678 640266 445774 640282
rect 445900 640714 446300 641094
rect 446397 641526 446493 641542
rect 446397 640982 446413 641526
rect 446477 640982 446493 641526
rect 446397 640966 446493 640982
rect 446620 641414 447020 641794
rect 447116 642226 447212 642242
rect 447116 641682 447132 642226
rect 447196 641682 447212 642226
rect 447116 641666 447212 641682
rect 447340 642114 447740 642494
rect 447835 642926 447931 642942
rect 447835 642382 447851 642926
rect 447915 642382 447931 642926
rect 447835 642366 447931 642382
rect 448060 642814 448460 643194
rect 448554 643626 448650 643642
rect 448554 643082 448570 643626
rect 448634 643082 448650 643626
rect 448554 643066 448650 643082
rect 448780 643514 449180 643894
rect 449273 643782 449289 644326
rect 449353 643782 449369 644326
rect 449992 644326 450088 644342
rect 449273 643766 449369 643782
rect 449500 644214 449900 644254
rect 449500 643894 449533 644214
rect 449853 643894 449900 644214
rect 448780 643194 448814 643514
rect 449134 643194 449180 643514
rect 448060 642494 448095 642814
rect 448415 642494 448460 642814
rect 447340 641794 447376 642114
rect 447696 641794 447740 642114
rect 446620 641094 446657 641414
rect 446977 641094 447020 641414
rect 445900 640394 445938 640714
rect 446258 640394 446300 640714
rect 445180 639694 445219 640014
rect 445539 639694 445580 640014
rect 444460 638994 444500 639314
rect 444820 638994 444860 639314
rect 444460 638614 444860 638994
rect 444959 639426 445055 639442
rect 444959 638882 444975 639426
rect 445039 638882 445055 639426
rect 444959 638866 445055 638882
rect 445180 639314 445580 639694
rect 445678 640126 445774 640142
rect 445678 639582 445694 640126
rect 445758 639582 445774 640126
rect 445678 639566 445774 639582
rect 445900 640014 446300 640394
rect 446397 640826 446493 640842
rect 446397 640282 446413 640826
rect 446477 640282 446493 640826
rect 446397 640266 446493 640282
rect 446620 640714 447020 641094
rect 447116 641526 447212 641542
rect 447116 640982 447132 641526
rect 447196 640982 447212 641526
rect 447116 640966 447212 640982
rect 447340 641414 447740 641794
rect 447835 642226 447931 642242
rect 447835 641682 447851 642226
rect 447915 641682 447931 642226
rect 447835 641666 447931 641682
rect 448060 642114 448460 642494
rect 448554 642926 448650 642942
rect 448554 642382 448570 642926
rect 448634 642382 448650 642926
rect 448554 642366 448650 642382
rect 448780 642814 449180 643194
rect 449273 643626 449369 643642
rect 449273 643082 449289 643626
rect 449353 643082 449369 643626
rect 449273 643066 449369 643082
rect 449500 643514 449900 643894
rect 449992 643782 450008 644326
rect 450072 643782 450088 644326
rect 450711 644326 450807 644342
rect 449992 643766 450088 643782
rect 450220 644214 450620 644254
rect 450220 643894 450252 644214
rect 450572 643894 450620 644214
rect 449500 643194 449533 643514
rect 449853 643194 449900 643514
rect 448780 642494 448814 642814
rect 449134 642494 449180 642814
rect 448060 641794 448095 642114
rect 448415 641794 448460 642114
rect 447340 641094 447376 641414
rect 447696 641094 447740 641414
rect 446620 640394 446657 640714
rect 446977 640394 447020 640714
rect 445900 639694 445938 640014
rect 446258 639694 446300 640014
rect 445180 638994 445219 639314
rect 445539 638994 445580 639314
rect 422960 638358 439052 638422
rect 422960 638294 437900 638358
rect 437964 638294 438028 638358
rect 438092 638294 438156 638358
rect 438220 638294 438284 638358
rect 438348 638294 438412 638358
rect 438476 638294 438540 638358
rect 438604 638294 438668 638358
rect 438732 638294 438796 638358
rect 438860 638294 438924 638358
rect 438988 638294 439052 638358
rect 422960 638230 439052 638294
rect 422960 638166 437900 638230
rect 437964 638166 438028 638230
rect 438092 638166 438156 638230
rect 438220 638166 438284 638230
rect 438348 638166 438412 638230
rect 438476 638166 438540 638230
rect 438604 638166 438668 638230
rect 438732 638166 438796 638230
rect 438860 638166 438924 638230
rect 438988 638166 439052 638230
rect 422960 638102 439052 638166
rect 422960 638038 437900 638102
rect 437964 638038 438028 638102
rect 438092 638038 438156 638102
rect 438220 638038 438284 638102
rect 438348 638038 438412 638102
rect 438476 638038 438540 638102
rect 438604 638038 438668 638102
rect 438732 638038 438796 638102
rect 438860 638038 438924 638102
rect 438988 638038 439052 638102
rect 422960 637974 439052 638038
rect 422960 637910 437900 637974
rect 437964 637910 438028 637974
rect 438092 637910 438156 637974
rect 438220 637910 438284 637974
rect 438348 637910 438412 637974
rect 438476 637910 438540 637974
rect 438604 637910 438668 637974
rect 438732 637910 438796 637974
rect 438860 637910 438924 637974
rect 438988 637910 439052 637974
rect 422960 637846 439052 637910
rect 444460 638294 444500 638614
rect 444820 638294 444860 638614
rect 444460 637914 444860 638294
rect 444959 638726 445055 638742
rect 444959 638182 444975 638726
rect 445039 638182 445055 638726
rect 444959 638166 445055 638182
rect 445180 638614 445580 638994
rect 445678 639426 445774 639442
rect 445678 638882 445694 639426
rect 445758 638882 445774 639426
rect 445678 638866 445774 638882
rect 445900 639314 446300 639694
rect 446397 640126 446493 640142
rect 446397 639582 446413 640126
rect 446477 639582 446493 640126
rect 446397 639566 446493 639582
rect 446620 640014 447020 640394
rect 447116 640826 447212 640842
rect 447116 640282 447132 640826
rect 447196 640282 447212 640826
rect 447116 640266 447212 640282
rect 447340 640714 447740 641094
rect 447835 641526 447931 641542
rect 447835 640982 447851 641526
rect 447915 640982 447931 641526
rect 447835 640966 447931 640982
rect 448060 641414 448460 641794
rect 448554 642226 448650 642242
rect 448554 641682 448570 642226
rect 448634 641682 448650 642226
rect 448554 641666 448650 641682
rect 448780 642114 449180 642494
rect 449273 642926 449369 642942
rect 449273 642382 449289 642926
rect 449353 642382 449369 642926
rect 449273 642366 449369 642382
rect 449500 642814 449900 643194
rect 449992 643626 450088 643642
rect 449992 643082 450008 643626
rect 450072 643082 450088 643626
rect 449992 643066 450088 643082
rect 450220 643514 450620 643894
rect 450711 643782 450727 644326
rect 450791 643782 450807 644326
rect 451430 644326 451526 644342
rect 450931 644214 451340 644254
rect 450931 643894 450971 644214
rect 451291 643894 451340 644214
rect 450931 643854 451340 643894
rect 450711 643766 450807 643782
rect 450220 643194 450252 643514
rect 450572 643194 450620 643514
rect 449500 642494 449533 642814
rect 449853 642494 449900 642814
rect 448780 641794 448814 642114
rect 449134 641794 449180 642114
rect 448060 641094 448095 641414
rect 448415 641094 448460 641414
rect 447340 640394 447376 640714
rect 447696 640394 447740 640714
rect 446620 639694 446657 640014
rect 446977 639694 447020 640014
rect 445900 638994 445938 639314
rect 446258 638994 446300 639314
rect 445180 638294 445219 638614
rect 445539 638294 445580 638614
rect 444460 637594 444500 637914
rect 444820 637594 444860 637914
rect 444460 637386 444860 637594
rect 444959 638026 445055 638042
rect 444959 637482 444975 638026
rect 445039 637482 445055 638026
rect 444959 637466 445055 637482
rect 445180 637914 445580 638294
rect 445678 638726 445774 638742
rect 445678 638182 445694 638726
rect 445758 638182 445774 638726
rect 445678 638166 445774 638182
rect 445900 638614 446300 638994
rect 446397 639426 446493 639442
rect 446397 638882 446413 639426
rect 446477 638882 446493 639426
rect 446397 638866 446493 638882
rect 446620 639314 447020 639694
rect 447116 640126 447212 640142
rect 447116 639582 447132 640126
rect 447196 639582 447212 640126
rect 447116 639566 447212 639582
rect 447340 640014 447740 640394
rect 447835 640826 447931 640842
rect 447835 640282 447851 640826
rect 447915 640282 447931 640826
rect 447835 640266 447931 640282
rect 448060 640714 448460 641094
rect 448554 641526 448650 641542
rect 448554 640982 448570 641526
rect 448634 640982 448650 641526
rect 448554 640966 448650 640982
rect 448780 641414 449180 641794
rect 449273 642226 449369 642242
rect 449273 641682 449289 642226
rect 449353 641682 449369 642226
rect 449273 641666 449369 641682
rect 449500 642114 449900 642494
rect 449992 642926 450088 642942
rect 449992 642382 450008 642926
rect 450072 642382 450088 642926
rect 449992 642366 450088 642382
rect 450220 642814 450620 643194
rect 450711 643626 450807 643642
rect 450711 643082 450727 643626
rect 450791 643082 450807 643626
rect 450711 643066 450807 643082
rect 450940 643514 451340 643854
rect 451430 643782 451446 644326
rect 451510 643782 451526 644326
rect 451430 643766 451526 643782
rect 482038 644254 482174 644354
rect 482274 644254 482398 644354
rect 482498 644254 482622 644354
rect 482722 644254 482846 644354
rect 482946 644254 483070 644354
rect 483170 644254 487200 644354
rect 482038 644130 487200 644254
rect 482038 644030 482174 644130
rect 482274 644030 482398 644130
rect 482498 644030 482622 644130
rect 482722 644030 482846 644130
rect 482946 644030 483070 644130
rect 483170 644030 487200 644130
rect 482038 644000 487200 644030
rect 491984 644000 492674 649744
rect 482038 643906 492674 644000
rect 482038 643806 482174 643906
rect 482274 643806 482398 643906
rect 482498 643806 482622 643906
rect 482722 643806 482846 643906
rect 482946 643806 483070 643906
rect 483170 643806 492674 643906
rect 482038 643682 492674 643806
rect 450940 643194 450971 643514
rect 451291 643194 451340 643514
rect 450220 642494 450252 642814
rect 450572 642494 450620 642814
rect 449500 641794 449533 642114
rect 449853 641794 449900 642114
rect 448780 641094 448814 641414
rect 449134 641094 449180 641414
rect 448060 640394 448095 640714
rect 448415 640394 448460 640714
rect 447340 639694 447376 640014
rect 447696 639694 447740 640014
rect 446620 638994 446657 639314
rect 446977 638994 447020 639314
rect 445900 638294 445938 638614
rect 446258 638294 446300 638614
rect 445180 637594 445219 637914
rect 445539 637594 445580 637914
rect 445180 637386 445580 637594
rect 445678 638026 445774 638042
rect 445678 637482 445694 638026
rect 445758 637482 445774 638026
rect 445678 637466 445774 637482
rect 445900 637914 446300 638294
rect 446397 638726 446493 638742
rect 446397 638182 446413 638726
rect 446477 638182 446493 638726
rect 446397 638166 446493 638182
rect 446620 638614 447020 638994
rect 447116 639426 447212 639442
rect 447116 638882 447132 639426
rect 447196 638882 447212 639426
rect 447116 638866 447212 638882
rect 447340 639314 447740 639694
rect 447835 640126 447931 640142
rect 447835 639582 447851 640126
rect 447915 639582 447931 640126
rect 447835 639566 447931 639582
rect 448060 640014 448460 640394
rect 448554 640826 448650 640842
rect 448554 640282 448570 640826
rect 448634 640282 448650 640826
rect 448554 640266 448650 640282
rect 448780 640714 449180 641094
rect 449273 641526 449369 641542
rect 449273 640982 449289 641526
rect 449353 640982 449369 641526
rect 449273 640966 449369 640982
rect 449500 641414 449900 641794
rect 449992 642226 450088 642242
rect 449992 641682 450008 642226
rect 450072 641682 450088 642226
rect 449992 641666 450088 641682
rect 450220 642114 450620 642494
rect 450711 642926 450807 642942
rect 450711 642382 450727 642926
rect 450791 642382 450807 642926
rect 450711 642366 450807 642382
rect 450940 642814 451340 643194
rect 451430 643626 451526 643642
rect 451430 643082 451446 643626
rect 451510 643082 451526 643626
rect 482038 643582 482174 643682
rect 482274 643582 482398 643682
rect 482498 643582 482622 643682
rect 482722 643582 482846 643682
rect 482946 643582 483070 643682
rect 483170 643582 492674 643682
rect 482038 643526 492674 643582
rect 451430 643066 451526 643082
rect 450940 642494 450971 642814
rect 451291 642494 451340 642814
rect 450220 641794 450252 642114
rect 450572 641794 450620 642114
rect 449500 641094 449533 641414
rect 449853 641094 449900 641414
rect 448780 640394 448814 640714
rect 449134 640394 449180 640714
rect 448060 639694 448095 640014
rect 448415 639694 448460 640014
rect 447340 638994 447376 639314
rect 447696 638994 447740 639314
rect 446620 638294 446657 638614
rect 446977 638294 447020 638614
rect 445900 637594 445938 637914
rect 446258 637594 446300 637914
rect 445900 637386 446300 637594
rect 446397 638026 446493 638042
rect 446397 637482 446413 638026
rect 446477 637482 446493 638026
rect 446397 637466 446493 637482
rect 446620 637914 447020 638294
rect 447116 638726 447212 638742
rect 447116 638182 447132 638726
rect 447196 638182 447212 638726
rect 447116 638166 447212 638182
rect 447340 638614 447740 638994
rect 447835 639426 447931 639442
rect 447835 638882 447851 639426
rect 447915 638882 447931 639426
rect 447835 638866 447931 638882
rect 448060 639314 448460 639694
rect 448554 640126 448650 640142
rect 448554 639582 448570 640126
rect 448634 639582 448650 640126
rect 448554 639566 448650 639582
rect 448780 640014 449180 640394
rect 449273 640826 449369 640842
rect 449273 640282 449289 640826
rect 449353 640282 449369 640826
rect 449273 640266 449369 640282
rect 449500 640714 449900 641094
rect 449992 641526 450088 641542
rect 449992 640982 450008 641526
rect 450072 640982 450088 641526
rect 449992 640966 450088 640982
rect 450220 641414 450620 641794
rect 450711 642226 450807 642242
rect 450711 641682 450727 642226
rect 450791 641682 450807 642226
rect 450711 641666 450807 641682
rect 450940 642114 451340 642494
rect 451430 642926 451526 642942
rect 451430 642382 451446 642926
rect 451510 642382 451526 642926
rect 451430 642366 451526 642382
rect 450940 641794 450971 642114
rect 451291 641794 451340 642114
rect 450220 641094 450252 641414
rect 450572 641094 450620 641414
rect 449500 640394 449533 640714
rect 449853 640394 449900 640714
rect 448780 639694 448814 640014
rect 449134 639694 449180 640014
rect 448060 638994 448095 639314
rect 448415 638994 448460 639314
rect 447340 638294 447376 638614
rect 447696 638294 447740 638614
rect 446620 637594 446657 637914
rect 446977 637594 447020 637914
rect 446620 637386 447020 637594
rect 447116 638026 447212 638042
rect 447116 637482 447132 638026
rect 447196 637482 447212 638026
rect 447116 637466 447212 637482
rect 447340 637914 447740 638294
rect 447835 638726 447931 638742
rect 447835 638182 447851 638726
rect 447915 638182 447931 638726
rect 447835 638166 447931 638182
rect 448060 638614 448460 638994
rect 448554 639426 448650 639442
rect 448554 638882 448570 639426
rect 448634 638882 448650 639426
rect 448554 638866 448650 638882
rect 448780 639314 449180 639694
rect 449273 640126 449369 640142
rect 449273 639582 449289 640126
rect 449353 639582 449369 640126
rect 449273 639566 449369 639582
rect 449500 640014 449900 640394
rect 449992 640826 450088 640842
rect 449992 640282 450008 640826
rect 450072 640282 450088 640826
rect 449992 640266 450088 640282
rect 450220 640714 450620 641094
rect 450711 641526 450807 641542
rect 450711 640982 450727 641526
rect 450791 640982 450807 641526
rect 450711 640966 450807 640982
rect 450940 641414 451340 641794
rect 451430 642226 451526 642242
rect 451430 641682 451446 642226
rect 451510 641682 451526 642226
rect 451430 641666 451526 641682
rect 450940 641094 450971 641414
rect 451291 641094 451340 641414
rect 450220 640394 450252 640714
rect 450572 640394 450620 640714
rect 449500 639694 449533 640014
rect 449853 639694 449900 640014
rect 448780 638994 448814 639314
rect 449134 638994 449180 639314
rect 448060 638294 448095 638614
rect 448415 638294 448460 638614
rect 447340 637594 447376 637914
rect 447696 637594 447740 637914
rect 447340 637386 447740 637594
rect 447835 638026 447931 638042
rect 447835 637482 447851 638026
rect 447915 637482 447931 638026
rect 447835 637466 447931 637482
rect 448060 637914 448460 638294
rect 448554 638726 448650 638742
rect 448554 638182 448570 638726
rect 448634 638182 448650 638726
rect 448554 638166 448650 638182
rect 448780 638614 449180 638994
rect 449273 639426 449369 639442
rect 449273 638882 449289 639426
rect 449353 638882 449369 639426
rect 449273 638866 449369 638882
rect 449500 639314 449900 639694
rect 449992 640126 450088 640142
rect 449992 639582 450008 640126
rect 450072 639582 450088 640126
rect 449992 639566 450088 639582
rect 450220 640014 450620 640394
rect 450711 640826 450807 640842
rect 450711 640282 450727 640826
rect 450791 640282 450807 640826
rect 450711 640266 450807 640282
rect 450940 640714 451340 641094
rect 451430 641526 451526 641542
rect 451430 640982 451446 641526
rect 451510 640982 451526 641526
rect 451430 640966 451526 640982
rect 459443 641050 459645 641051
rect 459443 640850 459444 641050
rect 459644 640850 459645 641050
rect 459443 640849 459645 640850
rect 459877 641050 460079 641051
rect 459877 640850 459878 641050
rect 460078 640850 460079 641050
rect 459877 640849 460079 640850
rect 460311 641050 460513 641051
rect 460311 640850 460312 641050
rect 460512 640850 460513 641050
rect 460311 640849 460513 640850
rect 460745 641050 460947 641051
rect 460745 640850 460746 641050
rect 460946 640850 460947 641050
rect 460745 640849 460947 640850
rect 461179 641050 461381 641051
rect 461179 640850 461180 641050
rect 461380 640850 461381 641050
rect 461179 640849 461381 640850
rect 461613 641050 461815 641051
rect 461613 640850 461614 641050
rect 461814 640850 461815 641050
rect 461613 640849 461815 640850
rect 462047 641050 462249 641051
rect 462047 640850 462048 641050
rect 462248 640850 462249 641050
rect 462047 640849 462249 640850
rect 462481 641050 462683 641051
rect 462481 640850 462482 641050
rect 462682 640850 462683 641050
rect 462481 640849 462683 640850
rect 462915 641050 463117 641051
rect 462915 640850 462916 641050
rect 463116 640850 463117 641050
rect 462915 640849 463117 640850
rect 463349 641050 463551 641051
rect 463349 640850 463350 641050
rect 463550 640850 463551 641050
rect 463349 640849 463551 640850
rect 463783 641050 463985 641051
rect 463783 640850 463784 641050
rect 463984 640850 463985 641050
rect 463783 640849 463985 640850
rect 464183 641050 464385 641051
rect 464183 640850 464184 641050
rect 464384 640850 464385 641050
rect 464183 640849 464385 640850
rect 464583 641050 464785 641051
rect 464583 640850 464584 641050
rect 464784 640850 464785 641050
rect 464583 640849 464785 640850
rect 464983 641050 465185 641051
rect 464983 640850 464984 641050
rect 465184 640850 465185 641050
rect 464983 640849 465185 640850
rect 465383 641050 465585 641051
rect 465383 640850 465384 641050
rect 465584 640850 465585 641050
rect 465383 640849 465585 640850
rect 465783 641050 465985 641051
rect 465783 640850 465784 641050
rect 465984 640850 465985 641050
rect 465783 640849 465985 640850
rect 466183 641050 466385 641051
rect 466183 640850 466184 641050
rect 466384 640850 466385 641050
rect 466183 640849 466385 640850
rect 466583 641050 466785 641051
rect 466583 640850 466584 641050
rect 466784 640850 466785 641050
rect 466583 640849 466785 640850
rect 466983 641050 467185 641051
rect 466983 640850 466984 641050
rect 467184 640850 467185 641050
rect 466983 640849 467185 640850
rect 467383 641050 467585 641051
rect 467383 640850 467384 641050
rect 467584 640850 467585 641050
rect 467383 640849 467585 640850
rect 468983 641050 469185 641051
rect 468983 640850 468984 641050
rect 469184 640850 469185 641050
rect 468983 640849 469185 640850
rect 469383 641050 469585 641051
rect 469383 640850 469384 641050
rect 469584 640850 469585 641050
rect 469383 640849 469585 640850
rect 469783 641050 469985 641051
rect 469783 640850 469784 641050
rect 469984 640850 469985 641050
rect 469783 640849 469985 640850
rect 470183 641050 470385 641051
rect 470183 640850 470184 641050
rect 470384 640850 470385 641050
rect 470183 640849 470385 640850
rect 470583 641050 470785 641051
rect 470583 640850 470584 641050
rect 470784 640850 470785 641050
rect 470583 640849 470785 640850
rect 470983 641050 471185 641051
rect 470983 640850 470984 641050
rect 471184 640850 471185 641050
rect 470983 640849 471185 640850
rect 471383 641050 471585 641051
rect 471383 640850 471384 641050
rect 471584 640850 471585 641050
rect 471383 640849 471585 640850
rect 471783 641050 471985 641051
rect 471783 640850 471784 641050
rect 471984 640850 471985 641050
rect 471783 640849 471985 640850
rect 472183 641050 472385 641051
rect 472183 640850 472184 641050
rect 472384 640850 472385 641050
rect 472183 640849 472385 640850
rect 450940 640394 450971 640714
rect 451291 640394 451340 640714
rect 450220 639694 450252 640014
rect 450572 639694 450620 640014
rect 449500 638994 449533 639314
rect 449853 638994 449900 639314
rect 448780 638294 448814 638614
rect 449134 638294 449180 638614
rect 448060 637594 448095 637914
rect 448415 637594 448460 637914
rect 448060 637386 448460 637594
rect 448554 638026 448650 638042
rect 448554 637482 448570 638026
rect 448634 637482 448650 638026
rect 448554 637466 448650 637482
rect 448780 637914 449180 638294
rect 449273 638726 449369 638742
rect 449273 638182 449289 638726
rect 449353 638182 449369 638726
rect 449273 638166 449369 638182
rect 449500 638614 449900 638994
rect 449992 639426 450088 639442
rect 449992 638882 450008 639426
rect 450072 638882 450088 639426
rect 449992 638866 450088 638882
rect 450220 639314 450620 639694
rect 450711 640126 450807 640142
rect 450711 639582 450727 640126
rect 450791 639582 450807 640126
rect 450711 639566 450807 639582
rect 450940 640014 451340 640394
rect 451430 640826 451526 640842
rect 451430 640282 451446 640826
rect 451510 640282 451526 640826
rect 459443 640616 459645 640617
rect 459443 640416 459444 640616
rect 459644 640416 459645 640616
rect 459443 640415 459645 640416
rect 459877 640616 460079 640617
rect 459877 640416 459878 640616
rect 460078 640416 460079 640616
rect 459877 640415 460079 640416
rect 460311 640616 460513 640617
rect 460311 640416 460312 640616
rect 460512 640416 460513 640616
rect 460311 640415 460513 640416
rect 460745 640616 460947 640617
rect 460745 640416 460746 640616
rect 460946 640416 460947 640616
rect 460745 640415 460947 640416
rect 461179 640616 461381 640617
rect 461179 640416 461180 640616
rect 461380 640416 461381 640616
rect 461179 640415 461381 640416
rect 461613 640616 461815 640617
rect 461613 640416 461614 640616
rect 461814 640416 461815 640616
rect 461613 640415 461815 640416
rect 462047 640616 462249 640617
rect 462047 640416 462048 640616
rect 462248 640416 462249 640616
rect 462047 640415 462249 640416
rect 462481 640616 462683 640617
rect 462481 640416 462482 640616
rect 462682 640416 462683 640616
rect 462481 640415 462683 640416
rect 462915 640616 463117 640617
rect 462915 640416 462916 640616
rect 463116 640416 463117 640616
rect 462915 640415 463117 640416
rect 463349 640616 463551 640617
rect 463349 640416 463350 640616
rect 463550 640416 463551 640616
rect 463349 640415 463551 640416
rect 463783 640616 463985 640617
rect 463783 640416 463784 640616
rect 463984 640416 463985 640616
rect 463783 640415 463985 640416
rect 451430 640266 451526 640282
rect 459443 640182 459645 640183
rect 450940 639694 450971 640014
rect 451291 639694 451340 640014
rect 450220 638994 450252 639314
rect 450572 638994 450620 639314
rect 449500 638294 449533 638614
rect 449853 638294 449900 638614
rect 448780 637594 448814 637914
rect 449134 637594 449180 637914
rect 448780 637386 449180 637594
rect 449273 638026 449369 638042
rect 449273 637482 449289 638026
rect 449353 637482 449369 638026
rect 449273 637466 449369 637482
rect 449500 637914 449900 638294
rect 449992 638726 450088 638742
rect 449992 638182 450008 638726
rect 450072 638182 450088 638726
rect 449992 638166 450088 638182
rect 450220 638614 450620 638994
rect 450711 639426 450807 639442
rect 450711 638882 450727 639426
rect 450791 638882 450807 639426
rect 450711 638866 450807 638882
rect 450940 639314 451340 639694
rect 451430 640126 451526 640142
rect 451430 639582 451446 640126
rect 451510 639582 451526 640126
rect 459443 639982 459444 640182
rect 459644 639982 459645 640182
rect 459443 639981 459645 639982
rect 459877 640182 460079 640183
rect 459877 639982 459878 640182
rect 460078 639982 460079 640182
rect 459877 639981 460079 639982
rect 460311 640182 460513 640183
rect 460311 639982 460312 640182
rect 460512 639982 460513 640182
rect 460311 639981 460513 639982
rect 460745 640182 460947 640183
rect 460745 639982 460746 640182
rect 460946 639982 460947 640182
rect 460745 639981 460947 639982
rect 461179 640182 461381 640183
rect 461179 639982 461180 640182
rect 461380 639982 461381 640182
rect 461179 639981 461381 639982
rect 461613 640182 461815 640183
rect 461613 639982 461614 640182
rect 461814 639982 461815 640182
rect 461613 639981 461815 639982
rect 462047 640182 462249 640183
rect 462047 639982 462048 640182
rect 462248 639982 462249 640182
rect 462047 639981 462249 639982
rect 462481 640182 462683 640183
rect 462481 639982 462482 640182
rect 462682 639982 462683 640182
rect 462481 639981 462683 639982
rect 462915 640182 463117 640183
rect 462915 639982 462916 640182
rect 463116 639982 463117 640182
rect 462915 639981 463117 639982
rect 463349 640182 463551 640183
rect 463349 639982 463350 640182
rect 463550 639982 463551 640182
rect 463349 639981 463551 639982
rect 463783 640182 463985 640183
rect 463783 639982 463784 640182
rect 463984 639982 463985 640182
rect 463783 639981 463985 639982
rect 451430 639566 451526 639582
rect 453001 639468 473313 639469
rect 450940 638994 450971 639314
rect 451291 638994 451340 639314
rect 450220 638294 450252 638614
rect 450572 638294 450620 638614
rect 449500 637594 449533 637914
rect 449853 637594 449900 637914
rect 449500 637386 449900 637594
rect 449992 638026 450088 638042
rect 449992 637482 450008 638026
rect 450072 637482 450088 638026
rect 449992 637466 450088 637482
rect 450220 637914 450620 638294
rect 450711 638726 450807 638742
rect 450711 638182 450727 638726
rect 450791 638182 450807 638726
rect 450711 638166 450807 638182
rect 450940 638614 451340 638994
rect 451430 639426 451526 639442
rect 451430 638882 451446 639426
rect 451510 638882 451526 639426
rect 451430 638866 451526 638882
rect 450940 638294 450971 638614
rect 451291 638294 451340 638614
rect 450220 637594 450252 637914
rect 450572 637594 450620 637914
rect 450220 637386 450620 637594
rect 450711 638026 450807 638042
rect 450711 637482 450727 638026
rect 450791 637482 450807 638026
rect 450711 637466 450807 637482
rect 450940 637914 451340 638294
rect 451430 638726 451526 638742
rect 451430 638182 451446 638726
rect 451510 638182 451526 638726
rect 453001 638496 453002 639468
rect 473312 638496 473313 639468
rect 453001 638495 473313 638496
rect 451430 638166 451526 638182
rect 450940 637594 450971 637914
rect 451291 637594 451340 637914
rect 450940 637394 451340 637594
rect 451430 638026 451526 638042
rect 451430 637482 451446 638026
rect 451510 637482 451526 638026
rect 451430 637466 451526 637482
rect 450940 637386 451360 637394
rect 444460 637379 451360 637386
rect 429064 636778 438924 636802
rect 429064 636678 437894 636778
rect 437994 636678 438118 636778
rect 438218 636678 438342 636778
rect 438442 636678 438566 636778
rect 438666 636678 438790 636778
rect 438890 636678 438924 636778
rect 429064 636554 438924 636678
rect 429064 636454 437894 636554
rect 437994 636454 438118 636554
rect 438218 636454 438342 636554
rect 438442 636454 438566 636554
rect 438666 636454 438790 636554
rect 438890 636454 438924 636554
rect 429064 636330 438924 636454
rect 429064 636230 437894 636330
rect 437994 636230 438118 636330
rect 438218 636230 438342 636330
rect 438442 636230 438566 636330
rect 438666 636230 438790 636330
rect 438890 636230 438924 636330
rect 429064 636106 438924 636230
rect 429064 636006 437894 636106
rect 437994 636006 438118 636106
rect 438218 636006 438342 636106
rect 438442 636006 438566 636106
rect 438666 636006 438790 636106
rect 438890 636006 438924 636106
rect 429064 635966 438924 636006
rect 429064 630222 429964 635966
rect 434748 635882 438924 635966
rect 434748 635782 437894 635882
rect 437994 635782 438118 635882
rect 438218 635782 438342 635882
rect 438442 635782 438566 635882
rect 438666 635782 438790 635882
rect 438890 635782 438924 635882
rect 434748 635658 438924 635782
rect 434748 635558 437894 635658
rect 437994 635558 438118 635658
rect 438218 635558 438342 635658
rect 438442 635558 438566 635658
rect 438666 635558 438790 635658
rect 438890 635558 438924 635658
rect 434748 635434 438924 635558
rect 434748 635334 437894 635434
rect 437994 635334 438118 635434
rect 438218 635334 438342 635434
rect 438442 635334 438566 635434
rect 438666 635334 438790 635434
rect 438890 635334 438924 635434
rect 434748 635210 438924 635334
rect 434748 635110 437894 635210
rect 437994 635110 438118 635210
rect 438218 635110 438342 635210
rect 438442 635110 438566 635210
rect 438666 635110 438790 635210
rect 438890 635110 438924 635210
rect 434748 634986 438924 635110
rect 434748 634886 437894 634986
rect 437994 634886 438118 634986
rect 438218 634886 438342 634986
rect 438442 634886 438566 634986
rect 438666 634886 438790 634986
rect 438890 634886 438924 634986
rect 434748 634762 438924 634886
rect 434748 634662 437894 634762
rect 437994 634662 438118 634762
rect 438218 634662 438342 634762
rect 438442 634662 438566 634762
rect 438666 634662 438790 634762
rect 438890 634662 438924 634762
rect 434748 634538 438924 634662
rect 434748 634438 437894 634538
rect 437994 634438 438118 634538
rect 438218 634438 438342 634538
rect 438442 634438 438566 634538
rect 438666 634438 438790 634538
rect 438890 634438 438924 634538
rect 434748 634314 438924 634438
rect 434748 634214 437894 634314
rect 437994 634214 438118 634314
rect 438218 634214 438342 634314
rect 438442 634214 438566 634314
rect 438666 634214 438790 634314
rect 438890 634214 438924 634314
rect 434748 634090 438924 634214
rect 434748 633990 437894 634090
rect 437994 633990 438118 634090
rect 438218 633990 438342 634090
rect 438442 633990 438566 634090
rect 438666 633990 438790 634090
rect 438890 633990 438924 634090
rect 434748 633866 438924 633990
rect 434748 633766 437894 633866
rect 437994 633766 438118 633866
rect 438218 633766 438342 633866
rect 438442 633766 438566 633866
rect 438666 633766 438790 633866
rect 438890 633766 438924 633866
rect 434748 633642 438924 633766
rect 434748 633542 437894 633642
rect 437994 633542 438118 633642
rect 438218 633542 438342 633642
rect 438442 633542 438566 633642
rect 438666 633542 438790 633642
rect 438890 633542 438924 633642
rect 434748 633418 438924 633542
rect 434748 633318 437894 633418
rect 437994 633318 438118 633418
rect 438218 633318 438342 633418
rect 438442 633318 438566 633418
rect 438666 633318 438790 633418
rect 438890 633318 438924 633418
rect 434748 633194 438924 633318
rect 434748 633094 437894 633194
rect 437994 633094 438118 633194
rect 438218 633094 438342 633194
rect 438442 633094 438566 633194
rect 438666 633094 438790 633194
rect 438890 633094 438924 633194
rect 434748 632970 438924 633094
rect 434748 632870 437894 632970
rect 437994 632870 438118 632970
rect 438218 632870 438342 632970
rect 438442 632870 438566 632970
rect 438666 632870 438790 632970
rect 438890 632870 438924 632970
rect 434748 632746 438924 632870
rect 434748 632646 437894 632746
rect 437994 632646 438118 632746
rect 438218 632646 438342 632746
rect 438442 632646 438566 632746
rect 438666 632646 438790 632746
rect 438890 632646 438924 632746
rect 434748 632522 438924 632646
rect 434748 632422 437894 632522
rect 437994 632422 438118 632522
rect 438218 632422 438342 632522
rect 438442 632422 438566 632522
rect 438666 632422 438790 632522
rect 438890 632422 438924 632522
rect 434748 632298 438924 632422
rect 443634 632333 452766 637379
rect 434748 632198 437894 632298
rect 437994 632198 438118 632298
rect 438218 632198 438342 632298
rect 438442 632198 438566 632298
rect 438666 632198 438790 632298
rect 438890 632198 438924 632298
rect 434748 632074 438924 632198
rect 434748 631974 437894 632074
rect 437994 631974 438118 632074
rect 438218 631974 438342 632074
rect 438442 631974 438566 632074
rect 438666 631974 438790 632074
rect 438890 631974 438924 632074
rect 443632 632331 452766 632333
rect 443632 632051 443634 632331
rect 444262 632051 452125 632331
rect 452753 632051 452766 632331
rect 443632 632049 452766 632051
rect 443634 632048 452766 632049
rect 482044 636778 492674 636788
rect 482044 636678 482174 636778
rect 482274 636678 482398 636778
rect 482498 636678 482622 636778
rect 482722 636678 482846 636778
rect 482946 636678 483070 636778
rect 483170 636678 492674 636778
rect 482044 636554 492674 636678
rect 482044 636454 482174 636554
rect 482274 636454 482398 636554
rect 482498 636454 482622 636554
rect 482722 636454 482846 636554
rect 482946 636454 483070 636554
rect 483170 636454 492674 636554
rect 482044 636344 492674 636454
rect 482044 636330 487200 636344
rect 482044 636230 482174 636330
rect 482274 636230 482398 636330
rect 482498 636230 482622 636330
rect 482722 636230 482846 636330
rect 482946 636230 483070 636330
rect 483170 636230 487200 636330
rect 482044 636106 487200 636230
rect 482044 636006 482174 636106
rect 482274 636006 482398 636106
rect 482498 636006 482622 636106
rect 482722 636006 482846 636106
rect 482946 636006 483070 636106
rect 483170 636006 487200 636106
rect 482044 635882 487200 636006
rect 482044 635782 482174 635882
rect 482274 635782 482398 635882
rect 482498 635782 482622 635882
rect 482722 635782 482846 635882
rect 482946 635782 483070 635882
rect 483170 635782 487200 635882
rect 482044 635658 487200 635782
rect 482044 635558 482174 635658
rect 482274 635558 482398 635658
rect 482498 635558 482622 635658
rect 482722 635558 482846 635658
rect 482946 635558 483070 635658
rect 483170 635558 487200 635658
rect 482044 635434 487200 635558
rect 482044 635334 482174 635434
rect 482274 635334 482398 635434
rect 482498 635334 482622 635434
rect 482722 635334 482846 635434
rect 482946 635334 483070 635434
rect 483170 635334 487200 635434
rect 482044 635210 487200 635334
rect 482044 635110 482174 635210
rect 482274 635110 482398 635210
rect 482498 635110 482622 635210
rect 482722 635110 482846 635210
rect 482946 635110 483070 635210
rect 483170 635110 487200 635210
rect 482044 634986 487200 635110
rect 482044 634886 482174 634986
rect 482274 634886 482398 634986
rect 482498 634886 482622 634986
rect 482722 634886 482846 634986
rect 482946 634886 483070 634986
rect 483170 634886 487200 634986
rect 482044 634762 487200 634886
rect 482044 634662 482174 634762
rect 482274 634662 482398 634762
rect 482498 634662 482622 634762
rect 482722 634662 482846 634762
rect 482946 634662 483070 634762
rect 483170 634662 487200 634762
rect 482044 634538 487200 634662
rect 482044 634438 482174 634538
rect 482274 634438 482398 634538
rect 482498 634438 482622 634538
rect 482722 634438 482846 634538
rect 482946 634438 483070 634538
rect 483170 634438 487200 634538
rect 482044 634314 487200 634438
rect 482044 634214 482174 634314
rect 482274 634214 482398 634314
rect 482498 634214 482622 634314
rect 482722 634214 482846 634314
rect 482946 634214 483070 634314
rect 483170 634214 487200 634314
rect 482044 634090 487200 634214
rect 482044 633990 482174 634090
rect 482274 633990 482398 634090
rect 482498 633990 482622 634090
rect 482722 633990 482846 634090
rect 482946 633990 483070 634090
rect 483170 633990 487200 634090
rect 482044 633866 487200 633990
rect 482044 633766 482174 633866
rect 482274 633766 482398 633866
rect 482498 633766 482622 633866
rect 482722 633766 482846 633866
rect 482946 633766 483070 633866
rect 483170 633766 487200 633866
rect 482044 633642 487200 633766
rect 482044 633542 482174 633642
rect 482274 633542 482398 633642
rect 482498 633542 482622 633642
rect 482722 633542 482846 633642
rect 482946 633542 483070 633642
rect 483170 633542 487200 633642
rect 482044 633418 487200 633542
rect 482044 633318 482174 633418
rect 482274 633318 482398 633418
rect 482498 633318 482622 633418
rect 482722 633318 482846 633418
rect 482946 633318 483070 633418
rect 483170 633318 487200 633418
rect 482044 633194 487200 633318
rect 482044 633094 482174 633194
rect 482274 633094 482398 633194
rect 482498 633094 482622 633194
rect 482722 633094 482846 633194
rect 482946 633094 483070 633194
rect 483170 633094 487200 633194
rect 482044 632970 487200 633094
rect 482044 632870 482174 632970
rect 482274 632870 482398 632970
rect 482498 632870 482622 632970
rect 482722 632870 482846 632970
rect 482946 632870 483070 632970
rect 483170 632870 487200 632970
rect 482044 632746 487200 632870
rect 482044 632646 482174 632746
rect 482274 632646 482398 632746
rect 482498 632646 482622 632746
rect 482722 632646 482846 632746
rect 482946 632646 483070 632746
rect 483170 632646 487200 632746
rect 482044 632522 487200 632646
rect 482044 632422 482174 632522
rect 482274 632422 482398 632522
rect 482498 632422 482622 632522
rect 482722 632422 482846 632522
rect 482946 632422 483070 632522
rect 483170 632422 487200 632522
rect 482044 632298 487200 632422
rect 482044 632198 482174 632298
rect 482274 632198 482398 632298
rect 482498 632198 482622 632298
rect 482722 632198 482846 632298
rect 482946 632198 483070 632298
rect 483170 632198 487200 632298
rect 482044 632074 487200 632198
rect 434748 631850 438924 631974
rect 434748 631750 437894 631850
rect 437994 631750 438118 631850
rect 438218 631750 438342 631850
rect 438442 631750 438566 631850
rect 438666 631750 438790 631850
rect 438890 631750 438924 631850
rect 434748 631626 438924 631750
rect 434748 631526 437894 631626
rect 437994 631526 438118 631626
rect 438218 631526 438342 631626
rect 438442 631526 438566 631626
rect 438666 631526 438790 631626
rect 438890 631526 438924 631626
rect 434748 631402 438924 631526
rect 434748 631302 437894 631402
rect 437994 631302 438118 631402
rect 438218 631302 438342 631402
rect 438442 631302 438566 631402
rect 438666 631302 438790 631402
rect 438890 631302 438924 631402
rect 434748 631178 438924 631302
rect 434748 631078 437894 631178
rect 437994 631078 438118 631178
rect 438218 631078 438342 631178
rect 438442 631078 438566 631178
rect 438666 631078 438790 631178
rect 438890 631078 438924 631178
rect 434748 630954 438924 631078
rect 434748 630854 437894 630954
rect 437994 630854 438118 630954
rect 438218 630854 438342 630954
rect 438442 630854 438566 630954
rect 438666 630854 438790 630954
rect 438890 630854 438924 630954
rect 434748 630730 438924 630854
rect 434748 630630 437894 630730
rect 437994 630630 438118 630730
rect 438218 630630 438342 630730
rect 438442 630630 438566 630730
rect 438666 630630 438790 630730
rect 438890 630630 438924 630730
rect 434748 630506 438924 630630
rect 434748 630406 437894 630506
rect 437994 630406 438118 630506
rect 438218 630406 438342 630506
rect 438442 630406 438566 630506
rect 438666 630406 438790 630506
rect 438890 630406 438924 630506
rect 434748 630282 438924 630406
rect 434748 630222 437894 630282
rect 429064 630182 437894 630222
rect 437994 630182 438118 630282
rect 438218 630182 438342 630282
rect 438442 630182 438566 630282
rect 438666 630182 438790 630282
rect 438890 630182 438924 630282
rect 429064 630122 438924 630182
rect 482044 631974 482174 632074
rect 482274 631974 482398 632074
rect 482498 631974 482622 632074
rect 482722 631974 482846 632074
rect 482946 631974 483070 632074
rect 483170 631974 487200 632074
rect 482044 631850 487200 631974
rect 482044 631750 482174 631850
rect 482274 631750 482398 631850
rect 482498 631750 482622 631850
rect 482722 631750 482846 631850
rect 482946 631750 483070 631850
rect 483170 631750 487200 631850
rect 482044 631626 487200 631750
rect 482044 631526 482174 631626
rect 482274 631526 482398 631626
rect 482498 631526 482622 631626
rect 482722 631526 482846 631626
rect 482946 631526 483070 631626
rect 483170 631526 487200 631626
rect 482044 631402 487200 631526
rect 482044 631302 482174 631402
rect 482274 631302 482398 631402
rect 482498 631302 482622 631402
rect 482722 631302 482846 631402
rect 482946 631302 483070 631402
rect 483170 631302 487200 631402
rect 482044 631178 487200 631302
rect 482044 631078 482174 631178
rect 482274 631078 482398 631178
rect 482498 631078 482622 631178
rect 482722 631078 482846 631178
rect 482946 631078 483070 631178
rect 483170 631078 487200 631178
rect 482044 630954 487200 631078
rect 482044 630854 482174 630954
rect 482274 630854 482398 630954
rect 482498 630854 482622 630954
rect 482722 630854 482846 630954
rect 482946 630854 483070 630954
rect 483170 630854 487200 630954
rect 482044 630730 487200 630854
rect 482044 630630 482174 630730
rect 482274 630630 482398 630730
rect 482498 630630 482622 630730
rect 482722 630630 482846 630730
rect 482946 630630 483070 630730
rect 483170 630630 487200 630730
rect 482044 630600 487200 630630
rect 491984 630600 492674 636344
rect 482044 630506 492674 630600
rect 482044 630406 482174 630506
rect 482274 630406 482398 630506
rect 482498 630406 482622 630506
rect 482722 630406 482846 630506
rect 482946 630406 483070 630506
rect 483170 630406 492674 630506
rect 482044 630282 492674 630406
rect 482044 630182 482174 630282
rect 482274 630182 482398 630282
rect 482498 630182 482622 630282
rect 482722 630182 482846 630282
rect 482946 630182 483070 630282
rect 483170 630182 492674 630282
rect 482044 630126 492674 630182
rect 475604 627681 482260 627686
rect 475604 627676 482261 627681
rect 438864 627661 445520 627666
rect 449334 627661 455990 627666
rect 438864 627656 445521 627661
rect 438864 627556 438920 627656
rect 439020 627556 439144 627656
rect 439244 627556 439368 627656
rect 439468 627556 439592 627656
rect 439692 627556 439816 627656
rect 439916 627556 440040 627656
rect 440140 627556 440264 627656
rect 440364 627556 440488 627656
rect 440588 627556 440712 627656
rect 440812 627556 440936 627656
rect 441036 627556 441160 627656
rect 441260 627556 441384 627656
rect 441484 627556 441608 627656
rect 441708 627556 441832 627656
rect 441932 627556 442056 627656
rect 442156 627556 442280 627656
rect 442380 627556 442504 627656
rect 442604 627556 442728 627656
rect 442828 627556 442952 627656
rect 443052 627556 443176 627656
rect 443276 627556 443400 627656
rect 443500 627556 443624 627656
rect 443724 627556 443848 627656
rect 443948 627556 444072 627656
rect 444172 627556 444296 627656
rect 444396 627556 444520 627656
rect 444620 627556 444744 627656
rect 444844 627556 444968 627656
rect 445068 627556 445192 627656
rect 445292 627556 445416 627656
rect 445516 627556 445521 627656
rect 438864 627551 445521 627556
rect 449334 627656 455991 627661
rect 449334 627556 449390 627656
rect 449490 627556 449614 627656
rect 449714 627556 449838 627656
rect 449938 627556 450062 627656
rect 450162 627556 450286 627656
rect 450386 627556 450510 627656
rect 450610 627556 450734 627656
rect 450834 627556 450958 627656
rect 451058 627556 451182 627656
rect 451282 627556 451406 627656
rect 451506 627556 451630 627656
rect 451730 627556 451854 627656
rect 451954 627556 452078 627656
rect 452178 627556 452302 627656
rect 452402 627556 452526 627656
rect 452626 627556 452750 627656
rect 452850 627556 452974 627656
rect 453074 627556 453198 627656
rect 453298 627556 453422 627656
rect 453522 627556 453646 627656
rect 453746 627556 453870 627656
rect 453970 627556 454094 627656
rect 454194 627556 454318 627656
rect 454418 627556 454542 627656
rect 454642 627556 454766 627656
rect 454866 627556 454990 627656
rect 455090 627556 455214 627656
rect 455314 627556 455438 627656
rect 455538 627556 455662 627656
rect 455762 627556 455886 627656
rect 455986 627556 455991 627656
rect 449334 627551 455991 627556
rect 475604 627576 475660 627676
rect 475760 627576 475884 627676
rect 475984 627576 476108 627676
rect 476208 627576 476332 627676
rect 476432 627576 476556 627676
rect 476656 627576 476780 627676
rect 476880 627576 477004 627676
rect 477104 627576 477228 627676
rect 477328 627576 477452 627676
rect 477552 627576 477676 627676
rect 477776 627576 477900 627676
rect 478000 627576 478124 627676
rect 478224 627576 478348 627676
rect 478448 627576 478572 627676
rect 478672 627576 478796 627676
rect 478896 627576 479020 627676
rect 479120 627576 479244 627676
rect 479344 627576 479468 627676
rect 479568 627576 479692 627676
rect 479792 627576 479916 627676
rect 480016 627576 480140 627676
rect 480240 627576 480364 627676
rect 480464 627576 480588 627676
rect 480688 627576 480812 627676
rect 480912 627576 481036 627676
rect 481136 627576 481260 627676
rect 481360 627576 481484 627676
rect 481584 627576 481708 627676
rect 481808 627576 481932 627676
rect 482032 627576 482156 627676
rect 482256 627576 482261 627676
rect 475604 627571 482261 627576
rect 438864 627437 445520 627551
rect 449334 627437 455990 627551
rect 475604 627457 482260 627571
rect 475604 627452 482261 627457
rect 438864 627432 445521 627437
rect 438864 627332 438920 627432
rect 439020 627332 439144 627432
rect 439244 627332 439368 627432
rect 439468 627332 439592 627432
rect 439692 627332 439816 627432
rect 439916 627332 440040 627432
rect 440140 627332 440264 627432
rect 440364 627332 440488 627432
rect 440588 627332 440712 627432
rect 440812 627332 440936 627432
rect 441036 627332 441160 627432
rect 441260 627332 441384 627432
rect 441484 627332 441608 627432
rect 441708 627332 441832 627432
rect 441932 627332 442056 627432
rect 442156 627332 442280 627432
rect 442380 627332 442504 627432
rect 442604 627332 442728 627432
rect 442828 627332 442952 627432
rect 443052 627332 443176 627432
rect 443276 627332 443400 627432
rect 443500 627332 443624 627432
rect 443724 627332 443848 627432
rect 443948 627332 444072 627432
rect 444172 627332 444296 627432
rect 444396 627332 444520 627432
rect 444620 627332 444744 627432
rect 444844 627332 444968 627432
rect 445068 627332 445192 627432
rect 445292 627332 445416 627432
rect 445516 627332 445521 627432
rect 438864 627327 445521 627332
rect 449334 627432 455991 627437
rect 449334 627332 449390 627432
rect 449490 627332 449614 627432
rect 449714 627332 449838 627432
rect 449938 627332 450062 627432
rect 450162 627332 450286 627432
rect 450386 627332 450510 627432
rect 450610 627332 450734 627432
rect 450834 627332 450958 627432
rect 451058 627332 451182 627432
rect 451282 627332 451406 627432
rect 451506 627332 451630 627432
rect 451730 627332 451854 627432
rect 451954 627332 452078 627432
rect 452178 627332 452302 627432
rect 452402 627332 452526 627432
rect 452626 627332 452750 627432
rect 452850 627332 452974 627432
rect 453074 627332 453198 627432
rect 453298 627332 453422 627432
rect 453522 627332 453646 627432
rect 453746 627332 453870 627432
rect 453970 627332 454094 627432
rect 454194 627332 454318 627432
rect 454418 627332 454542 627432
rect 454642 627332 454766 627432
rect 454866 627332 454990 627432
rect 455090 627332 455214 627432
rect 455314 627332 455438 627432
rect 455538 627332 455662 627432
rect 455762 627332 455886 627432
rect 455986 627332 455991 627432
rect 449334 627327 455991 627332
rect 475604 627352 475660 627452
rect 475760 627352 475884 627452
rect 475984 627352 476108 627452
rect 476208 627352 476332 627452
rect 476432 627352 476556 627452
rect 476656 627352 476780 627452
rect 476880 627352 477004 627452
rect 477104 627352 477228 627452
rect 477328 627352 477452 627452
rect 477552 627352 477676 627452
rect 477776 627352 477900 627452
rect 478000 627352 478124 627452
rect 478224 627352 478348 627452
rect 478448 627352 478572 627452
rect 478672 627352 478796 627452
rect 478896 627352 479020 627452
rect 479120 627352 479244 627452
rect 479344 627352 479468 627452
rect 479568 627352 479692 627452
rect 479792 627352 479916 627452
rect 480016 627352 480140 627452
rect 480240 627352 480364 627452
rect 480464 627352 480588 627452
rect 480688 627352 480812 627452
rect 480912 627352 481036 627452
rect 481136 627352 481260 627452
rect 481360 627352 481484 627452
rect 481584 627352 481708 627452
rect 481808 627352 481932 627452
rect 482032 627352 482156 627452
rect 482256 627352 482261 627452
rect 475604 627347 482261 627352
rect 438864 627213 445520 627327
rect 449334 627213 455990 627327
rect 475604 627233 482260 627347
rect 475604 627228 482261 627233
rect 438864 627208 445521 627213
rect 438864 627108 438920 627208
rect 439020 627108 439144 627208
rect 439244 627108 439368 627208
rect 439468 627108 439592 627208
rect 439692 627108 439816 627208
rect 439916 627108 440040 627208
rect 440140 627108 440264 627208
rect 440364 627108 440488 627208
rect 440588 627108 440712 627208
rect 440812 627108 440936 627208
rect 441036 627108 441160 627208
rect 441260 627108 441384 627208
rect 441484 627108 441608 627208
rect 441708 627108 441832 627208
rect 441932 627108 442056 627208
rect 442156 627108 442280 627208
rect 442380 627108 442504 627208
rect 442604 627108 442728 627208
rect 442828 627108 442952 627208
rect 443052 627108 443176 627208
rect 443276 627108 443400 627208
rect 443500 627108 443624 627208
rect 443724 627108 443848 627208
rect 443948 627108 444072 627208
rect 444172 627108 444296 627208
rect 444396 627108 444520 627208
rect 444620 627108 444744 627208
rect 444844 627108 444968 627208
rect 445068 627108 445192 627208
rect 445292 627108 445416 627208
rect 445516 627108 445521 627208
rect 438864 627103 445521 627108
rect 449334 627208 455991 627213
rect 449334 627108 449390 627208
rect 449490 627108 449614 627208
rect 449714 627108 449838 627208
rect 449938 627108 450062 627208
rect 450162 627108 450286 627208
rect 450386 627108 450510 627208
rect 450610 627108 450734 627208
rect 450834 627108 450958 627208
rect 451058 627108 451182 627208
rect 451282 627108 451406 627208
rect 451506 627108 451630 627208
rect 451730 627108 451854 627208
rect 451954 627108 452078 627208
rect 452178 627108 452302 627208
rect 452402 627108 452526 627208
rect 452626 627108 452750 627208
rect 452850 627108 452974 627208
rect 453074 627108 453198 627208
rect 453298 627108 453422 627208
rect 453522 627108 453646 627208
rect 453746 627108 453870 627208
rect 453970 627108 454094 627208
rect 454194 627108 454318 627208
rect 454418 627108 454542 627208
rect 454642 627108 454766 627208
rect 454866 627108 454990 627208
rect 455090 627108 455214 627208
rect 455314 627108 455438 627208
rect 455538 627108 455662 627208
rect 455762 627108 455886 627208
rect 455986 627108 455991 627208
rect 449334 627103 455991 627108
rect 475604 627128 475660 627228
rect 475760 627128 475884 627228
rect 475984 627128 476108 627228
rect 476208 627128 476332 627228
rect 476432 627128 476556 627228
rect 476656 627128 476780 627228
rect 476880 627128 477004 627228
rect 477104 627128 477228 627228
rect 477328 627128 477452 627228
rect 477552 627128 477676 627228
rect 477776 627128 477900 627228
rect 478000 627128 478124 627228
rect 478224 627128 478348 627228
rect 478448 627128 478572 627228
rect 478672 627128 478796 627228
rect 478896 627128 479020 627228
rect 479120 627128 479244 627228
rect 479344 627128 479468 627228
rect 479568 627128 479692 627228
rect 479792 627128 479916 627228
rect 480016 627128 480140 627228
rect 480240 627128 480364 627228
rect 480464 627128 480588 627228
rect 480688 627128 480812 627228
rect 480912 627128 481036 627228
rect 481136 627128 481260 627228
rect 481360 627128 481484 627228
rect 481584 627128 481708 627228
rect 481808 627128 481932 627228
rect 482032 627128 482156 627228
rect 482256 627128 482261 627228
rect 475604 627123 482261 627128
rect 438864 626989 445520 627103
rect 449334 626989 455990 627103
rect 475604 627009 482260 627123
rect 475604 627004 482261 627009
rect 438864 626984 445521 626989
rect 438864 626884 438920 626984
rect 439020 626884 439144 626984
rect 439244 626884 439368 626984
rect 439468 626884 439592 626984
rect 439692 626884 439816 626984
rect 439916 626884 440040 626984
rect 440140 626884 440264 626984
rect 440364 626884 440488 626984
rect 440588 626884 440712 626984
rect 440812 626884 440936 626984
rect 441036 626884 441160 626984
rect 441260 626884 441384 626984
rect 441484 626884 441608 626984
rect 441708 626884 441832 626984
rect 441932 626884 442056 626984
rect 442156 626884 442280 626984
rect 442380 626884 442504 626984
rect 442604 626884 442728 626984
rect 442828 626884 442952 626984
rect 443052 626884 443176 626984
rect 443276 626884 443400 626984
rect 443500 626884 443624 626984
rect 443724 626884 443848 626984
rect 443948 626884 444072 626984
rect 444172 626884 444296 626984
rect 444396 626884 444520 626984
rect 444620 626884 444744 626984
rect 444844 626884 444968 626984
rect 445068 626884 445192 626984
rect 445292 626884 445416 626984
rect 445516 626884 445521 626984
rect 438864 626879 445521 626884
rect 449334 626984 455991 626989
rect 449334 626884 449390 626984
rect 449490 626884 449614 626984
rect 449714 626884 449838 626984
rect 449938 626884 450062 626984
rect 450162 626884 450286 626984
rect 450386 626884 450510 626984
rect 450610 626884 450734 626984
rect 450834 626884 450958 626984
rect 451058 626884 451182 626984
rect 451282 626884 451406 626984
rect 451506 626884 451630 626984
rect 451730 626884 451854 626984
rect 451954 626884 452078 626984
rect 452178 626884 452302 626984
rect 452402 626884 452526 626984
rect 452626 626884 452750 626984
rect 452850 626884 452974 626984
rect 453074 626884 453198 626984
rect 453298 626884 453422 626984
rect 453522 626884 453646 626984
rect 453746 626884 453870 626984
rect 453970 626884 454094 626984
rect 454194 626884 454318 626984
rect 454418 626884 454542 626984
rect 454642 626884 454766 626984
rect 454866 626884 454990 626984
rect 455090 626884 455214 626984
rect 455314 626884 455438 626984
rect 455538 626884 455662 626984
rect 455762 626884 455886 626984
rect 455986 626884 455991 626984
rect 449334 626879 455991 626884
rect 475604 626904 475660 627004
rect 475760 626904 475884 627004
rect 475984 626904 476108 627004
rect 476208 626904 476332 627004
rect 476432 626904 476556 627004
rect 476656 626904 476780 627004
rect 476880 626904 477004 627004
rect 477104 626904 477228 627004
rect 477328 626904 477452 627004
rect 477552 626904 477676 627004
rect 477776 626904 477900 627004
rect 478000 626904 478124 627004
rect 478224 626904 478348 627004
rect 478448 626904 478572 627004
rect 478672 626904 478796 627004
rect 478896 626904 479020 627004
rect 479120 626904 479244 627004
rect 479344 626904 479468 627004
rect 479568 626904 479692 627004
rect 479792 626904 479916 627004
rect 480016 626904 480140 627004
rect 480240 626904 480364 627004
rect 480464 626904 480588 627004
rect 480688 626904 480812 627004
rect 480912 626904 481036 627004
rect 481136 626904 481260 627004
rect 481360 626904 481484 627004
rect 481584 626904 481708 627004
rect 481808 626904 481932 627004
rect 482032 626904 482156 627004
rect 482256 626904 482261 627004
rect 475604 626899 482261 626904
rect 438864 626765 445520 626879
rect 449334 626765 455990 626879
rect 475604 626785 482260 626899
rect 475604 626780 482261 626785
rect 438864 626760 445521 626765
rect 438864 626660 438920 626760
rect 439020 626660 439144 626760
rect 439244 626660 439368 626760
rect 439468 626660 439592 626760
rect 439692 626660 439816 626760
rect 439916 626660 440040 626760
rect 440140 626660 440264 626760
rect 440364 626660 440488 626760
rect 440588 626660 440712 626760
rect 440812 626660 440936 626760
rect 441036 626660 441160 626760
rect 441260 626660 441384 626760
rect 441484 626660 441608 626760
rect 441708 626660 441832 626760
rect 441932 626660 442056 626760
rect 442156 626660 442280 626760
rect 442380 626660 442504 626760
rect 442604 626660 442728 626760
rect 442828 626660 442952 626760
rect 443052 626660 443176 626760
rect 443276 626660 443400 626760
rect 443500 626660 443624 626760
rect 443724 626660 443848 626760
rect 443948 626660 444072 626760
rect 444172 626660 444296 626760
rect 444396 626660 444520 626760
rect 444620 626660 444744 626760
rect 444844 626660 444968 626760
rect 445068 626660 445192 626760
rect 445292 626660 445416 626760
rect 445516 626660 445521 626760
rect 438864 626655 445521 626660
rect 449334 626760 455991 626765
rect 449334 626660 449390 626760
rect 449490 626660 449614 626760
rect 449714 626660 449838 626760
rect 449938 626660 450062 626760
rect 450162 626660 450286 626760
rect 450386 626660 450510 626760
rect 450610 626660 450734 626760
rect 450834 626660 450958 626760
rect 451058 626660 451182 626760
rect 451282 626660 451406 626760
rect 451506 626660 451630 626760
rect 451730 626660 451854 626760
rect 451954 626660 452078 626760
rect 452178 626660 452302 626760
rect 452402 626660 452526 626760
rect 452626 626660 452750 626760
rect 452850 626660 452974 626760
rect 453074 626660 453198 626760
rect 453298 626660 453422 626760
rect 453522 626660 453646 626760
rect 453746 626660 453870 626760
rect 453970 626660 454094 626760
rect 454194 626660 454318 626760
rect 454418 626660 454542 626760
rect 454642 626660 454766 626760
rect 454866 626660 454990 626760
rect 455090 626660 455214 626760
rect 455314 626660 455438 626760
rect 455538 626660 455662 626760
rect 455762 626660 455886 626760
rect 455986 626660 455991 626760
rect 449334 626655 455991 626660
rect 475604 626680 475660 626780
rect 475760 626680 475884 626780
rect 475984 626680 476108 626780
rect 476208 626680 476332 626780
rect 476432 626680 476556 626780
rect 476656 626680 476780 626780
rect 476880 626680 477004 626780
rect 477104 626680 477228 626780
rect 477328 626680 477452 626780
rect 477552 626680 477676 626780
rect 477776 626680 477900 626780
rect 478000 626680 478124 626780
rect 478224 626680 478348 626780
rect 478448 626680 478572 626780
rect 478672 626680 478796 626780
rect 478896 626680 479020 626780
rect 479120 626680 479244 626780
rect 479344 626680 479468 626780
rect 479568 626680 479692 626780
rect 479792 626680 479916 626780
rect 480016 626680 480140 626780
rect 480240 626680 480364 626780
rect 480464 626680 480588 626780
rect 480688 626680 480812 626780
rect 480912 626680 481036 626780
rect 481136 626680 481260 626780
rect 481360 626680 481484 626780
rect 481584 626680 481708 626780
rect 481808 626680 481932 626780
rect 482032 626680 482156 626780
rect 482256 626680 482261 626780
rect 475604 626675 482261 626680
rect 438864 626626 445520 626655
rect 449334 626626 455990 626655
rect 475604 626646 482260 626675
rect 456344 623358 502000 623388
rect 425844 623266 502000 623358
rect 425844 623262 476524 623266
rect 425844 622946 438964 623262
rect 425844 617202 429964 622946
rect 434748 617518 438964 622946
rect 443748 617518 444964 623262
rect 449748 617518 450964 623262
rect 455748 617522 476524 623262
rect 481308 623144 502000 623266
rect 481308 617522 487200 623144
rect 455748 617518 487200 617522
rect 434748 617400 487200 617518
rect 491984 617400 502000 623144
rect 434748 617202 502000 617400
rect 425844 616726 502000 617202
rect 425844 616702 456344 616726
rect 456108 609506 502000 609988
rect 456108 603762 457524 609506
rect 462308 603762 465524 609506
rect 470308 603762 502000 609506
rect 456108 603422 502000 603762
rect 456104 603322 502000 603422
<< via4 >>
rect 453002 638496 473312 639468
<< mimcap2 >>
rect 440770 651454 441170 651494
rect 440770 651134 440810 651454
rect 441130 651134 441170 651454
rect 440770 651094 441170 651134
rect 441892 651454 442292 651494
rect 441892 651134 441932 651454
rect 442252 651134 442292 651454
rect 441892 651094 442292 651134
rect 443014 651454 443414 651494
rect 443014 651134 443054 651454
rect 443374 651134 443414 651454
rect 443014 651094 443414 651134
rect 444136 651454 444536 651494
rect 444136 651134 444176 651454
rect 444496 651134 444536 651454
rect 444136 651094 444536 651134
rect 445258 651454 445658 651494
rect 445258 651134 445298 651454
rect 445618 651134 445658 651454
rect 445258 651094 445658 651134
rect 446380 651454 446780 651494
rect 446380 651134 446420 651454
rect 446740 651134 446780 651454
rect 446380 651094 446780 651134
rect 447502 651454 447902 651494
rect 447502 651134 447542 651454
rect 447862 651134 447902 651454
rect 447502 651094 447902 651134
rect 448624 651454 449024 651494
rect 448624 651134 448664 651454
rect 448984 651134 449024 651454
rect 448624 651094 449024 651134
rect 449746 651454 450146 651494
rect 449746 651134 449786 651454
rect 450106 651134 450146 651454
rect 449746 651094 450146 651134
rect 450868 651454 451268 651494
rect 450868 651134 450908 651454
rect 451228 651134 451268 651454
rect 450868 651094 451268 651134
rect 440770 650754 441170 650794
rect 440770 650434 440810 650754
rect 441130 650434 441170 650754
rect 440770 650394 441170 650434
rect 441892 650754 442292 650794
rect 441892 650434 441932 650754
rect 442252 650434 442292 650754
rect 441892 650394 442292 650434
rect 443014 650754 443414 650794
rect 443014 650434 443054 650754
rect 443374 650434 443414 650754
rect 443014 650394 443414 650434
rect 444136 650754 444536 650794
rect 444136 650434 444176 650754
rect 444496 650434 444536 650754
rect 444136 650394 444536 650434
rect 445258 650754 445658 650794
rect 445258 650434 445298 650754
rect 445618 650434 445658 650754
rect 445258 650394 445658 650434
rect 446380 650754 446780 650794
rect 446380 650434 446420 650754
rect 446740 650434 446780 650754
rect 446380 650394 446780 650434
rect 447502 650754 447902 650794
rect 447502 650434 447542 650754
rect 447862 650434 447902 650754
rect 447502 650394 447902 650434
rect 448624 650754 449024 650794
rect 448624 650434 448664 650754
rect 448984 650434 449024 650754
rect 448624 650394 449024 650434
rect 449746 650754 450146 650794
rect 449746 650434 449786 650754
rect 450106 650434 450146 650754
rect 449746 650394 450146 650434
rect 450868 650754 451268 650794
rect 450868 650434 450908 650754
rect 451228 650434 451268 650754
rect 450868 650394 451268 650434
rect 440770 650054 441170 650094
rect 440770 649734 440810 650054
rect 441130 649734 441170 650054
rect 440770 649694 441170 649734
rect 441892 650054 442292 650094
rect 441892 649734 441932 650054
rect 442252 649734 442292 650054
rect 441892 649694 442292 649734
rect 443014 650054 443414 650094
rect 443014 649734 443054 650054
rect 443374 649734 443414 650054
rect 443014 649694 443414 649734
rect 444136 650054 444536 650094
rect 444136 649734 444176 650054
rect 444496 649734 444536 650054
rect 444136 649694 444536 649734
rect 445258 650054 445658 650094
rect 445258 649734 445298 650054
rect 445618 649734 445658 650054
rect 445258 649694 445658 649734
rect 446380 650054 446780 650094
rect 446380 649734 446420 650054
rect 446740 649734 446780 650054
rect 446380 649694 446780 649734
rect 447502 650054 447902 650094
rect 447502 649734 447542 650054
rect 447862 649734 447902 650054
rect 447502 649694 447902 649734
rect 448624 650054 449024 650094
rect 448624 649734 448664 650054
rect 448984 649734 449024 650054
rect 448624 649694 449024 649734
rect 449746 650054 450146 650094
rect 449746 649734 449786 650054
rect 450106 649734 450146 650054
rect 449746 649694 450146 649734
rect 450868 650054 451268 650094
rect 450868 649734 450908 650054
rect 451228 649734 451268 650054
rect 450868 649694 451268 649734
rect 440770 649354 441170 649394
rect 440770 649034 440810 649354
rect 441130 649034 441170 649354
rect 440770 648994 441170 649034
rect 441892 649354 442292 649394
rect 441892 649034 441932 649354
rect 442252 649034 442292 649354
rect 441892 648994 442292 649034
rect 443014 649354 443414 649394
rect 443014 649034 443054 649354
rect 443374 649034 443414 649354
rect 443014 648994 443414 649034
rect 444136 649354 444536 649394
rect 444136 649034 444176 649354
rect 444496 649034 444536 649354
rect 444136 648994 444536 649034
rect 445258 649354 445658 649394
rect 445258 649034 445298 649354
rect 445618 649034 445658 649354
rect 445258 648994 445658 649034
rect 446380 649354 446780 649394
rect 446380 649034 446420 649354
rect 446740 649034 446780 649354
rect 446380 648994 446780 649034
rect 447502 649354 447902 649394
rect 447502 649034 447542 649354
rect 447862 649034 447902 649354
rect 447502 648994 447902 649034
rect 448624 649354 449024 649394
rect 448624 649034 448664 649354
rect 448984 649034 449024 649354
rect 448624 648994 449024 649034
rect 449746 649354 450146 649394
rect 449746 649034 449786 649354
rect 450106 649034 450146 649354
rect 449746 648994 450146 649034
rect 450868 649354 451268 649394
rect 450868 649034 450908 649354
rect 451228 649034 451268 649354
rect 450868 648994 451268 649034
rect 440770 648654 441170 648694
rect 440770 648334 440810 648654
rect 441130 648334 441170 648654
rect 440770 648294 441170 648334
rect 441892 648654 442292 648694
rect 441892 648334 441932 648654
rect 442252 648334 442292 648654
rect 441892 648294 442292 648334
rect 443014 648654 443414 648694
rect 443014 648334 443054 648654
rect 443374 648334 443414 648654
rect 443014 648294 443414 648334
rect 444136 648654 444536 648694
rect 444136 648334 444176 648654
rect 444496 648334 444536 648654
rect 444136 648294 444536 648334
rect 445258 648654 445658 648694
rect 445258 648334 445298 648654
rect 445618 648334 445658 648654
rect 445258 648294 445658 648334
rect 446380 648654 446780 648694
rect 446380 648334 446420 648654
rect 446740 648334 446780 648654
rect 446380 648294 446780 648334
rect 447502 648654 447902 648694
rect 447502 648334 447542 648654
rect 447862 648334 447902 648654
rect 447502 648294 447902 648334
rect 448624 648654 449024 648694
rect 448624 648334 448664 648654
rect 448984 648334 449024 648654
rect 448624 648294 449024 648334
rect 449746 648654 450146 648694
rect 449746 648334 449786 648654
rect 450106 648334 450146 648654
rect 449746 648294 450146 648334
rect 450868 648654 451268 648694
rect 450868 648334 450908 648654
rect 451228 648334 451268 648654
rect 450868 648294 451268 648334
rect 440770 647954 441170 647994
rect 440770 647634 440810 647954
rect 441130 647634 441170 647954
rect 440770 647594 441170 647634
rect 441892 647954 442292 647994
rect 441892 647634 441932 647954
rect 442252 647634 442292 647954
rect 441892 647594 442292 647634
rect 443014 647954 443414 647994
rect 443014 647634 443054 647954
rect 443374 647634 443414 647954
rect 443014 647594 443414 647634
rect 444136 647954 444536 647994
rect 444136 647634 444176 647954
rect 444496 647634 444536 647954
rect 444136 647594 444536 647634
rect 445258 647954 445658 647994
rect 445258 647634 445298 647954
rect 445618 647634 445658 647954
rect 445258 647594 445658 647634
rect 446380 647954 446780 647994
rect 446380 647634 446420 647954
rect 446740 647634 446780 647954
rect 446380 647594 446780 647634
rect 447502 647954 447902 647994
rect 447502 647634 447542 647954
rect 447862 647634 447902 647954
rect 447502 647594 447902 647634
rect 448624 647954 449024 647994
rect 448624 647634 448664 647954
rect 448984 647634 449024 647954
rect 448624 647594 449024 647634
rect 449746 647954 450146 647994
rect 449746 647634 449786 647954
rect 450106 647634 450146 647954
rect 449746 647594 450146 647634
rect 450868 647954 451268 647994
rect 450868 647634 450908 647954
rect 451228 647634 451268 647954
rect 450868 647594 451268 647634
rect 440770 647254 441170 647294
rect 440770 646934 440810 647254
rect 441130 646934 441170 647254
rect 440770 646894 441170 646934
rect 441892 647254 442292 647294
rect 441892 646934 441932 647254
rect 442252 646934 442292 647254
rect 441892 646894 442292 646934
rect 443014 647254 443414 647294
rect 443014 646934 443054 647254
rect 443374 646934 443414 647254
rect 443014 646894 443414 646934
rect 444136 647254 444536 647294
rect 444136 646934 444176 647254
rect 444496 646934 444536 647254
rect 444136 646894 444536 646934
rect 445258 647254 445658 647294
rect 445258 646934 445298 647254
rect 445618 646934 445658 647254
rect 445258 646894 445658 646934
rect 446380 647254 446780 647294
rect 446380 646934 446420 647254
rect 446740 646934 446780 647254
rect 446380 646894 446780 646934
rect 447502 647254 447902 647294
rect 447502 646934 447542 647254
rect 447862 646934 447902 647254
rect 447502 646894 447902 646934
rect 448624 647254 449024 647294
rect 448624 646934 448664 647254
rect 448984 646934 449024 647254
rect 448624 646894 449024 646934
rect 449746 647254 450146 647294
rect 449746 646934 449786 647254
rect 450106 646934 450146 647254
rect 449746 646894 450146 646934
rect 450868 647254 451268 647294
rect 450868 646934 450908 647254
rect 451228 646934 451268 647254
rect 450868 646894 451268 646934
rect 440770 646554 441170 646594
rect 440770 646234 440810 646554
rect 441130 646234 441170 646554
rect 440770 646194 441170 646234
rect 441892 646554 442292 646594
rect 441892 646234 441932 646554
rect 442252 646234 442292 646554
rect 441892 646194 442292 646234
rect 443014 646554 443414 646594
rect 443014 646234 443054 646554
rect 443374 646234 443414 646554
rect 443014 646194 443414 646234
rect 444136 646554 444536 646594
rect 444136 646234 444176 646554
rect 444496 646234 444536 646554
rect 444136 646194 444536 646234
rect 445258 646554 445658 646594
rect 445258 646234 445298 646554
rect 445618 646234 445658 646554
rect 445258 646194 445658 646234
rect 446380 646554 446780 646594
rect 446380 646234 446420 646554
rect 446740 646234 446780 646554
rect 446380 646194 446780 646234
rect 447502 646554 447902 646594
rect 447502 646234 447542 646554
rect 447862 646234 447902 646554
rect 447502 646194 447902 646234
rect 448624 646554 449024 646594
rect 448624 646234 448664 646554
rect 448984 646234 449024 646554
rect 448624 646194 449024 646234
rect 449746 646554 450146 646594
rect 449746 646234 449786 646554
rect 450106 646234 450146 646554
rect 449746 646194 450146 646234
rect 450868 646554 451268 646594
rect 450868 646234 450908 646554
rect 451228 646234 451268 646554
rect 450868 646194 451268 646234
rect 440770 645854 441170 645894
rect 440770 645534 440810 645854
rect 441130 645534 441170 645854
rect 440770 645494 441170 645534
rect 441892 645854 442292 645894
rect 441892 645534 441932 645854
rect 442252 645534 442292 645854
rect 441892 645494 442292 645534
rect 443014 645854 443414 645894
rect 443014 645534 443054 645854
rect 443374 645534 443414 645854
rect 443014 645494 443414 645534
rect 444136 645854 444536 645894
rect 444136 645534 444176 645854
rect 444496 645534 444536 645854
rect 444136 645494 444536 645534
rect 445258 645854 445658 645894
rect 445258 645534 445298 645854
rect 445618 645534 445658 645854
rect 445258 645494 445658 645534
rect 446380 645854 446780 645894
rect 446380 645534 446420 645854
rect 446740 645534 446780 645854
rect 446380 645494 446780 645534
rect 447502 645854 447902 645894
rect 447502 645534 447542 645854
rect 447862 645534 447902 645854
rect 447502 645494 447902 645534
rect 448624 645854 449024 645894
rect 448624 645534 448664 645854
rect 448984 645534 449024 645854
rect 448624 645494 449024 645534
rect 449746 645854 450146 645894
rect 449746 645534 449786 645854
rect 450106 645534 450146 645854
rect 449746 645494 450146 645534
rect 450868 645854 451268 645894
rect 450868 645534 450908 645854
rect 451228 645534 451268 645854
rect 450868 645494 451268 645534
rect 440770 645154 441170 645194
rect 440770 644834 440810 645154
rect 441130 644834 441170 645154
rect 440770 644794 441170 644834
rect 441892 645154 442292 645194
rect 441892 644834 441932 645154
rect 442252 644834 442292 645154
rect 441892 644794 442292 644834
rect 443014 645154 443414 645194
rect 443014 644834 443054 645154
rect 443374 644834 443414 645154
rect 443014 644794 443414 644834
rect 444136 645154 444536 645194
rect 444136 644834 444176 645154
rect 444496 644834 444536 645154
rect 444136 644794 444536 644834
rect 445258 645154 445658 645194
rect 445258 644834 445298 645154
rect 445618 644834 445658 645154
rect 445258 644794 445658 644834
rect 446380 645154 446780 645194
rect 446380 644834 446420 645154
rect 446740 644834 446780 645154
rect 446380 644794 446780 644834
rect 447502 645154 447902 645194
rect 447502 644834 447542 645154
rect 447862 644834 447902 645154
rect 447502 644794 447902 644834
rect 448624 645154 449024 645194
rect 448624 644834 448664 645154
rect 448984 644834 449024 645154
rect 448624 644794 449024 644834
rect 449746 645154 450146 645194
rect 449746 644834 449786 645154
rect 450106 644834 450146 645154
rect 449746 644794 450146 644834
rect 450868 645154 451268 645194
rect 450868 644834 450908 645154
rect 451228 644834 451268 645154
rect 450868 644794 451268 644834
<< mimcap2contact >>
rect 440810 651134 441130 651454
rect 441932 651134 442252 651454
rect 443054 651134 443374 651454
rect 444176 651134 444496 651454
rect 445298 651134 445618 651454
rect 446420 651134 446740 651454
rect 447542 651134 447862 651454
rect 448664 651134 448984 651454
rect 449786 651134 450106 651454
rect 450908 651134 451228 651454
rect 440810 650434 441130 650754
rect 441932 650434 442252 650754
rect 443054 650434 443374 650754
rect 444176 650434 444496 650754
rect 445298 650434 445618 650754
rect 446420 650434 446740 650754
rect 447542 650434 447862 650754
rect 448664 650434 448984 650754
rect 449786 650434 450106 650754
rect 450908 650434 451228 650754
rect 440810 649734 441130 650054
rect 441932 649734 442252 650054
rect 443054 649734 443374 650054
rect 444176 649734 444496 650054
rect 445298 649734 445618 650054
rect 446420 649734 446740 650054
rect 447542 649734 447862 650054
rect 448664 649734 448984 650054
rect 449786 649734 450106 650054
rect 450908 649734 451228 650054
rect 440810 649034 441130 649354
rect 441932 649034 442252 649354
rect 443054 649034 443374 649354
rect 444176 649034 444496 649354
rect 445298 649034 445618 649354
rect 446420 649034 446740 649354
rect 447542 649034 447862 649354
rect 448664 649034 448984 649354
rect 449786 649034 450106 649354
rect 450908 649034 451228 649354
rect 440810 648334 441130 648654
rect 441932 648334 442252 648654
rect 443054 648334 443374 648654
rect 444176 648334 444496 648654
rect 445298 648334 445618 648654
rect 446420 648334 446740 648654
rect 447542 648334 447862 648654
rect 448664 648334 448984 648654
rect 449786 648334 450106 648654
rect 450908 648334 451228 648654
rect 440810 647634 441130 647954
rect 441932 647634 442252 647954
rect 443054 647634 443374 647954
rect 444176 647634 444496 647954
rect 445298 647634 445618 647954
rect 446420 647634 446740 647954
rect 447542 647634 447862 647954
rect 448664 647634 448984 647954
rect 449786 647634 450106 647954
rect 450908 647634 451228 647954
rect 440810 646934 441130 647254
rect 441932 646934 442252 647254
rect 443054 646934 443374 647254
rect 444176 646934 444496 647254
rect 445298 646934 445618 647254
rect 446420 646934 446740 647254
rect 447542 646934 447862 647254
rect 448664 646934 448984 647254
rect 449786 646934 450106 647254
rect 450908 646934 451228 647254
rect 440810 646234 441130 646554
rect 441932 646234 442252 646554
rect 443054 646234 443374 646554
rect 444176 646234 444496 646554
rect 445298 646234 445618 646554
rect 446420 646234 446740 646554
rect 447542 646234 447862 646554
rect 448664 646234 448984 646554
rect 449786 646234 450106 646554
rect 450908 646234 451228 646554
rect 440810 645534 441130 645854
rect 441932 645534 442252 645854
rect 443054 645534 443374 645854
rect 444176 645534 444496 645854
rect 445298 645534 445618 645854
rect 446420 645534 446740 645854
rect 447542 645534 447862 645854
rect 448664 645534 448984 645854
rect 449786 645534 450106 645854
rect 450908 645534 451228 645854
rect 440810 644834 441130 645154
rect 441932 644834 442252 645154
rect 443054 644834 443374 645154
rect 444176 644834 444496 645154
rect 445298 644834 445618 645154
rect 446420 644834 446740 645154
rect 447542 644834 447862 645154
rect 448664 644834 448984 645154
rect 449786 644834 450106 645154
rect 450908 644834 451228 645154
<< metal5 >>
rect 440716 651638 473330 651913
rect 440716 651454 473486 651638
rect 440716 651134 440810 651454
rect 441130 651134 441932 651454
rect 442252 651134 443054 651454
rect 443374 651134 444176 651454
rect 444496 651134 445298 651454
rect 445618 651134 446420 651454
rect 446740 651134 447542 651454
rect 447862 651134 448664 651454
rect 448984 651134 449786 651454
rect 450106 651134 450908 651454
rect 451228 651134 473486 651454
rect 440716 650754 473486 651134
rect 440716 650434 440810 650754
rect 441130 650434 441932 650754
rect 442252 650434 443054 650754
rect 443374 650434 444176 650754
rect 444496 650434 445298 650754
rect 445618 650434 446420 650754
rect 446740 650434 447542 650754
rect 447862 650434 448664 650754
rect 448984 650434 449786 650754
rect 450106 650434 450908 650754
rect 451228 650434 473486 650754
rect 440716 650054 473486 650434
rect 440716 649734 440810 650054
rect 441130 649734 441932 650054
rect 442252 649734 443054 650054
rect 443374 649734 444176 650054
rect 444496 649734 445298 650054
rect 445618 649734 446420 650054
rect 446740 649734 447542 650054
rect 447862 649734 448664 650054
rect 448984 649734 449786 650054
rect 450106 649734 450908 650054
rect 451228 649734 473486 650054
rect 440716 649354 473486 649734
rect 440716 649034 440810 649354
rect 441130 649034 441932 649354
rect 442252 649034 443054 649354
rect 443374 649034 444176 649354
rect 444496 649034 445298 649354
rect 445618 649034 446420 649354
rect 446740 649034 447542 649354
rect 447862 649034 448664 649354
rect 448984 649034 449786 649354
rect 450106 649034 450908 649354
rect 451228 649034 473486 649354
rect 440716 648654 473486 649034
rect 440716 648334 440810 648654
rect 441130 648334 441932 648654
rect 442252 648334 443054 648654
rect 443374 648334 444176 648654
rect 444496 648334 445298 648654
rect 445618 648334 446420 648654
rect 446740 648334 447542 648654
rect 447862 648334 448664 648654
rect 448984 648334 449786 648654
rect 450106 648334 450908 648654
rect 451228 648334 473486 648654
rect 440716 647954 473486 648334
rect 440716 647634 440810 647954
rect 441130 647634 441932 647954
rect 442252 647634 443054 647954
rect 443374 647634 444176 647954
rect 444496 647634 445298 647954
rect 445618 647634 446420 647954
rect 446740 647634 447542 647954
rect 447862 647634 448664 647954
rect 448984 647634 449786 647954
rect 450106 647634 450908 647954
rect 451228 647634 473486 647954
rect 440716 647254 473486 647634
rect 440716 646934 440810 647254
rect 441130 646934 441932 647254
rect 442252 646934 443054 647254
rect 443374 646934 444176 647254
rect 444496 646934 445298 647254
rect 445618 646934 446420 647254
rect 446740 646934 447542 647254
rect 447862 646934 448664 647254
rect 448984 646934 449786 647254
rect 450106 646934 450908 647254
rect 451228 646934 473486 647254
rect 440716 646554 473486 646934
rect 440716 646234 440810 646554
rect 441130 646234 441932 646554
rect 442252 646234 443054 646554
rect 443374 646234 444176 646554
rect 444496 646234 445298 646554
rect 445618 646234 446420 646554
rect 446740 646234 447542 646554
rect 447862 646234 448664 646554
rect 448984 646234 449786 646554
rect 450106 646234 450908 646554
rect 451228 646234 473486 646554
rect 440716 645854 473486 646234
rect 440716 645534 440810 645854
rect 441130 645534 441932 645854
rect 442252 645534 443054 645854
rect 443374 645534 444176 645854
rect 444496 645534 445298 645854
rect 445618 645534 446420 645854
rect 446740 645534 447542 645854
rect 447862 645534 448664 645854
rect 448984 645534 449786 645854
rect 450106 645534 450908 645854
rect 451228 645534 473486 645854
rect 440716 645154 473486 645534
rect 440716 644834 440810 645154
rect 441130 644834 441932 645154
rect 442252 644834 443054 645154
rect 443374 644834 444176 645154
rect 444496 644834 445298 645154
rect 445618 644834 446420 645154
rect 446740 644834 447542 645154
rect 447862 644834 448664 645154
rect 448984 644834 449786 645154
rect 450106 644834 450908 645154
rect 451228 644834 473486 645154
rect 440716 639468 473486 644834
rect 440716 638496 453002 639468
rect 473312 638496 473486 639468
rect 440716 638436 473486 638496
rect 453002 638398 473486 638436
<< res2p85 >>
rect 453314 644538 453888 647866
rect 454132 644538 454706 647866
rect 454950 644538 455524 647866
rect 456586 644948 457160 649252
rect 457404 644948 457978 649252
rect 458222 644948 458796 649252
rect 459040 644948 459614 649252
rect 461494 642882 462068 649190
rect 462312 642882 462886 649190
rect 463130 642882 463704 649190
rect 463948 642882 464522 649190
rect 464766 642882 465340 649190
rect 465584 642882 466158 649190
rect 466402 642882 466976 649190
rect 467220 642882 467794 649190
rect 468038 642882 468612 649190
rect 468856 642882 469430 649190
rect 469674 642882 470248 649190
rect 470492 642882 471066 649190
rect 471310 642882 471884 649190
rect 472128 642882 472702 649190
rect 472946 642882 473520 649190
rect 473764 642882 474338 649190
rect 474582 642882 475156 649190
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 7 1288
timestamp 1650294714
transform 1 0 474692 0 1 629606
box 0 0 1340 1340
<< labels >>
flabel metal1 442994 636190 443456 636388 1 FreeSans 1600 0 0 0 bandgaptop_flat_0/porst
flabel metal1 459390 640512 464058 641188 1 FreeSans 1600 0 0 0 bandgaptop_flat_0/Vbg
flabel metal2 440936 632416 442718 632486 1 FreeSans 800 0 0 0 bandgaptop_flat_0/ampcurrentsource_0/Vq
flabel metal2 440936 632626 442718 632696 1 FreeSans 800 0 0 0 bandgaptop_flat_0/ampcurrentsource_0/Vx
flabel locali 441796 633386 441878 633414 1 FreeSans 800 0 0 0 bandgaptop_flat_0/ampcurrentsource_0/GND!
flabel metal2 447688 629126 447704 629250 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/VDD!
flabel metal2 448342 632354 448358 632478 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vq
flabel metal2 448284 634614 448300 634694 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Va
flabel metal2 447512 634474 447528 634554 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vb
flabel metal2 449018 632058 449112 632324 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vgate
flabel metal2 447294 632058 447388 632324 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vgate
flabel metal1 445936 632072 445970 632164 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/vg
flabel metal2 450036 628926 450058 629050 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vx
flabel psubdiffcont 444814 632730 444914 634330 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/GND!
flabel psubdiff 450264 634330 450464 634430 5 FreeSans 800 180 0 0 bandgaptop_flat_0/amplifier_0/GND!
rlabel via1 454130 629106 454176 629150 5 bandgaptop_flat_0/currentmirror_0/Vgate
rlabel metal3 454852 628750 454986 628868 5 bandgaptop_flat_0/currentmirror_0/VDD!
flabel metal1 461658 637290 461958 637390 5 FreeSans 1600 0 0 0 bandgaptop_flat_0/currentmirror_0/Vbg
flabel metal2 461658 637890 461858 637990 5 FreeSans 1600 0 0 0 bandgaptop_flat_0/currentmirror_0/Vb
flabel via2 461658 638490 461858 638590 5 FreeSans 1600 0 0 0 bandgaptop_flat_0/currentmirror_0/Va
flabel metal2 463132 649188 463702 649620 1 FreeSans 800 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/VbEnd
flabel metal2 463950 642452 464520 642884 1 FreeSans 800 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/VbgEnd
flabel metal2 462314 648388 462884 649620 1 FreeSans 800 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/VaEnd
flabel metal2 472058 642186 472750 642878 1 FreeSans 1600 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/Vbg
flabel metal2 473688 642180 474392 642884 1 FreeSans 1600 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/Vb
flabel metal1 472870 641614 473574 642186 3 FreeSans 1600 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/Va
rlabel psubdiffcont 437892 626630 481132 627630 1 bandgaptop_flat_0/GND
rlabel metal3 441982 628688 442692 629110 1 bandgaptop_flat_0/VDD
flabel metal2 473854 629908 474990 630856 7 FreeSans 1600 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/Vbneg
<< end >>
