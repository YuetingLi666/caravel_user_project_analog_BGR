magic
tech sky130A
magscale 1 2
timestamp 1654929205
<< nwell >>
rect 575184 493285 580570 493663
rect 575183 492161 580570 493285
rect 574658 358981 580044 359359
rect 574657 357857 580044 358981
rect 575106 312813 580492 313191
rect 575105 311689 580492 312813
<< pwell >>
rect 560637 492423 565907 493475
rect 562136 492003 562308 492105
rect 563436 492003 563608 492105
rect 564736 492003 564908 492105
rect 565874 492003 565966 492175
rect 560573 403281 565843 404333
rect 562072 402861 562244 402963
rect 563372 402861 563544 402963
rect 564672 402861 564844 402963
rect 565810 402861 565902 403033
rect 560529 357963 565799 359015
rect 562028 357543 562200 357645
rect 563328 357543 563500 357645
rect 564628 357543 564800 357645
rect 565766 357543 565858 357715
rect 560391 311655 565661 312707
rect 561890 311235 562062 311337
rect 563190 311235 563362 311337
rect 564490 311235 564662 311337
rect 565628 311235 565720 311407
<< pmoslvt >>
rect 575277 492223 575477 493223
rect 575535 492223 575735 493223
rect 575793 492223 575993 493223
rect 576051 492223 576251 493223
rect 576309 492223 576509 493223
rect 576567 492223 576767 493223
rect 576825 492223 577025 493223
rect 577083 492223 577283 493223
rect 577341 492223 577541 493223
rect 577599 492223 577799 493223
rect 577857 492223 578057 493223
rect 578115 492223 578315 493223
rect 578373 492223 578573 493223
rect 578631 492223 578831 493223
rect 578889 492223 579089 493223
rect 579147 492223 579347 493223
rect 579405 492223 579605 493223
rect 579663 492223 579863 493223
rect 579921 492223 580121 493223
rect 580179 492223 580379 493223
rect 574751 357919 574951 358919
rect 575009 357919 575209 358919
rect 575267 357919 575467 358919
rect 575525 357919 575725 358919
rect 575783 357919 575983 358919
rect 576041 357919 576241 358919
rect 576299 357919 576499 358919
rect 576557 357919 576757 358919
rect 576815 357919 577015 358919
rect 577073 357919 577273 358919
rect 577331 357919 577531 358919
rect 577589 357919 577789 358919
rect 577847 357919 578047 358919
rect 578105 357919 578305 358919
rect 578363 357919 578563 358919
rect 578621 357919 578821 358919
rect 578879 357919 579079 358919
rect 579137 357919 579337 358919
rect 579395 357919 579595 358919
rect 579653 357919 579853 358919
rect 575199 311751 575399 312751
rect 575457 311751 575657 312751
rect 575715 311751 575915 312751
rect 575973 311751 576173 312751
rect 576231 311751 576431 312751
rect 576489 311751 576689 312751
rect 576747 311751 576947 312751
rect 577005 311751 577205 312751
rect 577263 311751 577463 312751
rect 577521 311751 577721 312751
rect 577779 311751 577979 312751
rect 578037 311751 578237 312751
rect 578295 311751 578495 312751
rect 578553 311751 578753 312751
rect 578811 311751 579011 312751
rect 579069 311751 579269 312751
rect 579327 311751 579527 312751
rect 579585 311751 579785 312751
rect 579843 311751 580043 312751
rect 580101 311751 580301 312751
<< nmoslvt >>
rect 560721 492449 560921 493449
rect 560979 492449 561179 493449
rect 561237 492449 561437 493449
rect 561495 492449 561695 493449
rect 561753 492449 561953 493449
rect 562011 492449 562211 493449
rect 562269 492449 562469 493449
rect 562527 492449 562727 493449
rect 562785 492449 562985 493449
rect 563043 492449 563243 493449
rect 563301 492449 563501 493449
rect 563559 492449 563759 493449
rect 563817 492449 564017 493449
rect 564075 492449 564275 493449
rect 564333 492449 564533 493449
rect 564591 492449 564791 493449
rect 564849 492449 565049 493449
rect 565107 492449 565307 493449
rect 565365 492449 565565 493449
rect 565623 492449 565823 493449
rect 560657 403307 560857 404307
rect 560915 403307 561115 404307
rect 561173 403307 561373 404307
rect 561431 403307 561631 404307
rect 561689 403307 561889 404307
rect 561947 403307 562147 404307
rect 562205 403307 562405 404307
rect 562463 403307 562663 404307
rect 562721 403307 562921 404307
rect 562979 403307 563179 404307
rect 563237 403307 563437 404307
rect 563495 403307 563695 404307
rect 563753 403307 563953 404307
rect 564011 403307 564211 404307
rect 564269 403307 564469 404307
rect 564527 403307 564727 404307
rect 564785 403307 564985 404307
rect 565043 403307 565243 404307
rect 565301 403307 565501 404307
rect 565559 403307 565759 404307
rect 560613 357989 560813 358989
rect 560871 357989 561071 358989
rect 561129 357989 561329 358989
rect 561387 357989 561587 358989
rect 561645 357989 561845 358989
rect 561903 357989 562103 358989
rect 562161 357989 562361 358989
rect 562419 357989 562619 358989
rect 562677 357989 562877 358989
rect 562935 357989 563135 358989
rect 563193 357989 563393 358989
rect 563451 357989 563651 358989
rect 563709 357989 563909 358989
rect 563967 357989 564167 358989
rect 564225 357989 564425 358989
rect 564483 357989 564683 358989
rect 564741 357989 564941 358989
rect 564999 357989 565199 358989
rect 565257 357989 565457 358989
rect 565515 357989 565715 358989
rect 560475 311681 560675 312681
rect 560733 311681 560933 312681
rect 560991 311681 561191 312681
rect 561249 311681 561449 312681
rect 561507 311681 561707 312681
rect 561765 311681 561965 312681
rect 562023 311681 562223 312681
rect 562281 311681 562481 312681
rect 562539 311681 562739 312681
rect 562797 311681 562997 312681
rect 563055 311681 563255 312681
rect 563313 311681 563513 312681
rect 563571 311681 563771 312681
rect 563829 311681 564029 312681
rect 564087 311681 564287 312681
rect 564345 311681 564545 312681
rect 564603 311681 564803 312681
rect 564861 311681 565061 312681
rect 565119 311681 565319 312681
rect 565377 311681 565577 312681
<< ndiff >>
rect 560663 493408 560721 493449
rect 560663 493374 560675 493408
rect 560709 493374 560721 493408
rect 560663 493340 560721 493374
rect 560663 493306 560675 493340
rect 560709 493306 560721 493340
rect 560663 493272 560721 493306
rect 560663 493238 560675 493272
rect 560709 493238 560721 493272
rect 560663 493204 560721 493238
rect 560663 493170 560675 493204
rect 560709 493170 560721 493204
rect 560663 493136 560721 493170
rect 560663 493102 560675 493136
rect 560709 493102 560721 493136
rect 560663 493068 560721 493102
rect 560663 493034 560675 493068
rect 560709 493034 560721 493068
rect 560663 493000 560721 493034
rect 560663 492966 560675 493000
rect 560709 492966 560721 493000
rect 560663 492932 560721 492966
rect 560663 492898 560675 492932
rect 560709 492898 560721 492932
rect 560663 492864 560721 492898
rect 560663 492830 560675 492864
rect 560709 492830 560721 492864
rect 560663 492796 560721 492830
rect 560663 492762 560675 492796
rect 560709 492762 560721 492796
rect 560663 492728 560721 492762
rect 560663 492694 560675 492728
rect 560709 492694 560721 492728
rect 560663 492660 560721 492694
rect 560663 492626 560675 492660
rect 560709 492626 560721 492660
rect 560663 492592 560721 492626
rect 560663 492558 560675 492592
rect 560709 492558 560721 492592
rect 560663 492524 560721 492558
rect 560663 492490 560675 492524
rect 560709 492490 560721 492524
rect 560663 492449 560721 492490
rect 560921 493408 560979 493449
rect 560921 493374 560933 493408
rect 560967 493374 560979 493408
rect 560921 493340 560979 493374
rect 560921 493306 560933 493340
rect 560967 493306 560979 493340
rect 560921 493272 560979 493306
rect 560921 493238 560933 493272
rect 560967 493238 560979 493272
rect 560921 493204 560979 493238
rect 560921 493170 560933 493204
rect 560967 493170 560979 493204
rect 560921 493136 560979 493170
rect 560921 493102 560933 493136
rect 560967 493102 560979 493136
rect 560921 493068 560979 493102
rect 560921 493034 560933 493068
rect 560967 493034 560979 493068
rect 560921 493000 560979 493034
rect 560921 492966 560933 493000
rect 560967 492966 560979 493000
rect 560921 492932 560979 492966
rect 560921 492898 560933 492932
rect 560967 492898 560979 492932
rect 560921 492864 560979 492898
rect 560921 492830 560933 492864
rect 560967 492830 560979 492864
rect 560921 492796 560979 492830
rect 560921 492762 560933 492796
rect 560967 492762 560979 492796
rect 560921 492728 560979 492762
rect 560921 492694 560933 492728
rect 560967 492694 560979 492728
rect 560921 492660 560979 492694
rect 560921 492626 560933 492660
rect 560967 492626 560979 492660
rect 560921 492592 560979 492626
rect 560921 492558 560933 492592
rect 560967 492558 560979 492592
rect 560921 492524 560979 492558
rect 560921 492490 560933 492524
rect 560967 492490 560979 492524
rect 560921 492449 560979 492490
rect 561179 493408 561237 493449
rect 561179 493374 561191 493408
rect 561225 493374 561237 493408
rect 561179 493340 561237 493374
rect 561179 493306 561191 493340
rect 561225 493306 561237 493340
rect 561179 493272 561237 493306
rect 561179 493238 561191 493272
rect 561225 493238 561237 493272
rect 561179 493204 561237 493238
rect 561179 493170 561191 493204
rect 561225 493170 561237 493204
rect 561179 493136 561237 493170
rect 561179 493102 561191 493136
rect 561225 493102 561237 493136
rect 561179 493068 561237 493102
rect 561179 493034 561191 493068
rect 561225 493034 561237 493068
rect 561179 493000 561237 493034
rect 561179 492966 561191 493000
rect 561225 492966 561237 493000
rect 561179 492932 561237 492966
rect 561179 492898 561191 492932
rect 561225 492898 561237 492932
rect 561179 492864 561237 492898
rect 561179 492830 561191 492864
rect 561225 492830 561237 492864
rect 561179 492796 561237 492830
rect 561179 492762 561191 492796
rect 561225 492762 561237 492796
rect 561179 492728 561237 492762
rect 561179 492694 561191 492728
rect 561225 492694 561237 492728
rect 561179 492660 561237 492694
rect 561179 492626 561191 492660
rect 561225 492626 561237 492660
rect 561179 492592 561237 492626
rect 561179 492558 561191 492592
rect 561225 492558 561237 492592
rect 561179 492524 561237 492558
rect 561179 492490 561191 492524
rect 561225 492490 561237 492524
rect 561179 492449 561237 492490
rect 561437 493408 561495 493449
rect 561437 493374 561449 493408
rect 561483 493374 561495 493408
rect 561437 493340 561495 493374
rect 561437 493306 561449 493340
rect 561483 493306 561495 493340
rect 561437 493272 561495 493306
rect 561437 493238 561449 493272
rect 561483 493238 561495 493272
rect 561437 493204 561495 493238
rect 561437 493170 561449 493204
rect 561483 493170 561495 493204
rect 561437 493136 561495 493170
rect 561437 493102 561449 493136
rect 561483 493102 561495 493136
rect 561437 493068 561495 493102
rect 561437 493034 561449 493068
rect 561483 493034 561495 493068
rect 561437 493000 561495 493034
rect 561437 492966 561449 493000
rect 561483 492966 561495 493000
rect 561437 492932 561495 492966
rect 561437 492898 561449 492932
rect 561483 492898 561495 492932
rect 561437 492864 561495 492898
rect 561437 492830 561449 492864
rect 561483 492830 561495 492864
rect 561437 492796 561495 492830
rect 561437 492762 561449 492796
rect 561483 492762 561495 492796
rect 561437 492728 561495 492762
rect 561437 492694 561449 492728
rect 561483 492694 561495 492728
rect 561437 492660 561495 492694
rect 561437 492626 561449 492660
rect 561483 492626 561495 492660
rect 561437 492592 561495 492626
rect 561437 492558 561449 492592
rect 561483 492558 561495 492592
rect 561437 492524 561495 492558
rect 561437 492490 561449 492524
rect 561483 492490 561495 492524
rect 561437 492449 561495 492490
rect 561695 493408 561753 493449
rect 561695 493374 561707 493408
rect 561741 493374 561753 493408
rect 561695 493340 561753 493374
rect 561695 493306 561707 493340
rect 561741 493306 561753 493340
rect 561695 493272 561753 493306
rect 561695 493238 561707 493272
rect 561741 493238 561753 493272
rect 561695 493204 561753 493238
rect 561695 493170 561707 493204
rect 561741 493170 561753 493204
rect 561695 493136 561753 493170
rect 561695 493102 561707 493136
rect 561741 493102 561753 493136
rect 561695 493068 561753 493102
rect 561695 493034 561707 493068
rect 561741 493034 561753 493068
rect 561695 493000 561753 493034
rect 561695 492966 561707 493000
rect 561741 492966 561753 493000
rect 561695 492932 561753 492966
rect 561695 492898 561707 492932
rect 561741 492898 561753 492932
rect 561695 492864 561753 492898
rect 561695 492830 561707 492864
rect 561741 492830 561753 492864
rect 561695 492796 561753 492830
rect 561695 492762 561707 492796
rect 561741 492762 561753 492796
rect 561695 492728 561753 492762
rect 561695 492694 561707 492728
rect 561741 492694 561753 492728
rect 561695 492660 561753 492694
rect 561695 492626 561707 492660
rect 561741 492626 561753 492660
rect 561695 492592 561753 492626
rect 561695 492558 561707 492592
rect 561741 492558 561753 492592
rect 561695 492524 561753 492558
rect 561695 492490 561707 492524
rect 561741 492490 561753 492524
rect 561695 492449 561753 492490
rect 561953 493408 562011 493449
rect 561953 493374 561965 493408
rect 561999 493374 562011 493408
rect 561953 493340 562011 493374
rect 561953 493306 561965 493340
rect 561999 493306 562011 493340
rect 561953 493272 562011 493306
rect 561953 493238 561965 493272
rect 561999 493238 562011 493272
rect 561953 493204 562011 493238
rect 561953 493170 561965 493204
rect 561999 493170 562011 493204
rect 561953 493136 562011 493170
rect 561953 493102 561965 493136
rect 561999 493102 562011 493136
rect 561953 493068 562011 493102
rect 561953 493034 561965 493068
rect 561999 493034 562011 493068
rect 561953 493000 562011 493034
rect 561953 492966 561965 493000
rect 561999 492966 562011 493000
rect 561953 492932 562011 492966
rect 561953 492898 561965 492932
rect 561999 492898 562011 492932
rect 561953 492864 562011 492898
rect 561953 492830 561965 492864
rect 561999 492830 562011 492864
rect 561953 492796 562011 492830
rect 561953 492762 561965 492796
rect 561999 492762 562011 492796
rect 561953 492728 562011 492762
rect 561953 492694 561965 492728
rect 561999 492694 562011 492728
rect 561953 492660 562011 492694
rect 561953 492626 561965 492660
rect 561999 492626 562011 492660
rect 561953 492592 562011 492626
rect 561953 492558 561965 492592
rect 561999 492558 562011 492592
rect 561953 492524 562011 492558
rect 561953 492490 561965 492524
rect 561999 492490 562011 492524
rect 561953 492449 562011 492490
rect 562211 493408 562269 493449
rect 562211 493374 562223 493408
rect 562257 493374 562269 493408
rect 562211 493340 562269 493374
rect 562211 493306 562223 493340
rect 562257 493306 562269 493340
rect 562211 493272 562269 493306
rect 562211 493238 562223 493272
rect 562257 493238 562269 493272
rect 562211 493204 562269 493238
rect 562211 493170 562223 493204
rect 562257 493170 562269 493204
rect 562211 493136 562269 493170
rect 562211 493102 562223 493136
rect 562257 493102 562269 493136
rect 562211 493068 562269 493102
rect 562211 493034 562223 493068
rect 562257 493034 562269 493068
rect 562211 493000 562269 493034
rect 562211 492966 562223 493000
rect 562257 492966 562269 493000
rect 562211 492932 562269 492966
rect 562211 492898 562223 492932
rect 562257 492898 562269 492932
rect 562211 492864 562269 492898
rect 562211 492830 562223 492864
rect 562257 492830 562269 492864
rect 562211 492796 562269 492830
rect 562211 492762 562223 492796
rect 562257 492762 562269 492796
rect 562211 492728 562269 492762
rect 562211 492694 562223 492728
rect 562257 492694 562269 492728
rect 562211 492660 562269 492694
rect 562211 492626 562223 492660
rect 562257 492626 562269 492660
rect 562211 492592 562269 492626
rect 562211 492558 562223 492592
rect 562257 492558 562269 492592
rect 562211 492524 562269 492558
rect 562211 492490 562223 492524
rect 562257 492490 562269 492524
rect 562211 492449 562269 492490
rect 562469 493408 562527 493449
rect 562469 493374 562481 493408
rect 562515 493374 562527 493408
rect 562469 493340 562527 493374
rect 562469 493306 562481 493340
rect 562515 493306 562527 493340
rect 562469 493272 562527 493306
rect 562469 493238 562481 493272
rect 562515 493238 562527 493272
rect 562469 493204 562527 493238
rect 562469 493170 562481 493204
rect 562515 493170 562527 493204
rect 562469 493136 562527 493170
rect 562469 493102 562481 493136
rect 562515 493102 562527 493136
rect 562469 493068 562527 493102
rect 562469 493034 562481 493068
rect 562515 493034 562527 493068
rect 562469 493000 562527 493034
rect 562469 492966 562481 493000
rect 562515 492966 562527 493000
rect 562469 492932 562527 492966
rect 562469 492898 562481 492932
rect 562515 492898 562527 492932
rect 562469 492864 562527 492898
rect 562469 492830 562481 492864
rect 562515 492830 562527 492864
rect 562469 492796 562527 492830
rect 562469 492762 562481 492796
rect 562515 492762 562527 492796
rect 562469 492728 562527 492762
rect 562469 492694 562481 492728
rect 562515 492694 562527 492728
rect 562469 492660 562527 492694
rect 562469 492626 562481 492660
rect 562515 492626 562527 492660
rect 562469 492592 562527 492626
rect 562469 492558 562481 492592
rect 562515 492558 562527 492592
rect 562469 492524 562527 492558
rect 562469 492490 562481 492524
rect 562515 492490 562527 492524
rect 562469 492449 562527 492490
rect 562727 493408 562785 493449
rect 562727 493374 562739 493408
rect 562773 493374 562785 493408
rect 562727 493340 562785 493374
rect 562727 493306 562739 493340
rect 562773 493306 562785 493340
rect 562727 493272 562785 493306
rect 562727 493238 562739 493272
rect 562773 493238 562785 493272
rect 562727 493204 562785 493238
rect 562727 493170 562739 493204
rect 562773 493170 562785 493204
rect 562727 493136 562785 493170
rect 562727 493102 562739 493136
rect 562773 493102 562785 493136
rect 562727 493068 562785 493102
rect 562727 493034 562739 493068
rect 562773 493034 562785 493068
rect 562727 493000 562785 493034
rect 562727 492966 562739 493000
rect 562773 492966 562785 493000
rect 562727 492932 562785 492966
rect 562727 492898 562739 492932
rect 562773 492898 562785 492932
rect 562727 492864 562785 492898
rect 562727 492830 562739 492864
rect 562773 492830 562785 492864
rect 562727 492796 562785 492830
rect 562727 492762 562739 492796
rect 562773 492762 562785 492796
rect 562727 492728 562785 492762
rect 562727 492694 562739 492728
rect 562773 492694 562785 492728
rect 562727 492660 562785 492694
rect 562727 492626 562739 492660
rect 562773 492626 562785 492660
rect 562727 492592 562785 492626
rect 562727 492558 562739 492592
rect 562773 492558 562785 492592
rect 562727 492524 562785 492558
rect 562727 492490 562739 492524
rect 562773 492490 562785 492524
rect 562727 492449 562785 492490
rect 562985 493408 563043 493449
rect 562985 493374 562997 493408
rect 563031 493374 563043 493408
rect 562985 493340 563043 493374
rect 562985 493306 562997 493340
rect 563031 493306 563043 493340
rect 562985 493272 563043 493306
rect 562985 493238 562997 493272
rect 563031 493238 563043 493272
rect 562985 493204 563043 493238
rect 562985 493170 562997 493204
rect 563031 493170 563043 493204
rect 562985 493136 563043 493170
rect 562985 493102 562997 493136
rect 563031 493102 563043 493136
rect 562985 493068 563043 493102
rect 562985 493034 562997 493068
rect 563031 493034 563043 493068
rect 562985 493000 563043 493034
rect 562985 492966 562997 493000
rect 563031 492966 563043 493000
rect 562985 492932 563043 492966
rect 562985 492898 562997 492932
rect 563031 492898 563043 492932
rect 562985 492864 563043 492898
rect 562985 492830 562997 492864
rect 563031 492830 563043 492864
rect 562985 492796 563043 492830
rect 562985 492762 562997 492796
rect 563031 492762 563043 492796
rect 562985 492728 563043 492762
rect 562985 492694 562997 492728
rect 563031 492694 563043 492728
rect 562985 492660 563043 492694
rect 562985 492626 562997 492660
rect 563031 492626 563043 492660
rect 562985 492592 563043 492626
rect 562985 492558 562997 492592
rect 563031 492558 563043 492592
rect 562985 492524 563043 492558
rect 562985 492490 562997 492524
rect 563031 492490 563043 492524
rect 562985 492449 563043 492490
rect 563243 493408 563301 493449
rect 563243 493374 563255 493408
rect 563289 493374 563301 493408
rect 563243 493340 563301 493374
rect 563243 493306 563255 493340
rect 563289 493306 563301 493340
rect 563243 493272 563301 493306
rect 563243 493238 563255 493272
rect 563289 493238 563301 493272
rect 563243 493204 563301 493238
rect 563243 493170 563255 493204
rect 563289 493170 563301 493204
rect 563243 493136 563301 493170
rect 563243 493102 563255 493136
rect 563289 493102 563301 493136
rect 563243 493068 563301 493102
rect 563243 493034 563255 493068
rect 563289 493034 563301 493068
rect 563243 493000 563301 493034
rect 563243 492966 563255 493000
rect 563289 492966 563301 493000
rect 563243 492932 563301 492966
rect 563243 492898 563255 492932
rect 563289 492898 563301 492932
rect 563243 492864 563301 492898
rect 563243 492830 563255 492864
rect 563289 492830 563301 492864
rect 563243 492796 563301 492830
rect 563243 492762 563255 492796
rect 563289 492762 563301 492796
rect 563243 492728 563301 492762
rect 563243 492694 563255 492728
rect 563289 492694 563301 492728
rect 563243 492660 563301 492694
rect 563243 492626 563255 492660
rect 563289 492626 563301 492660
rect 563243 492592 563301 492626
rect 563243 492558 563255 492592
rect 563289 492558 563301 492592
rect 563243 492524 563301 492558
rect 563243 492490 563255 492524
rect 563289 492490 563301 492524
rect 563243 492449 563301 492490
rect 563501 493408 563559 493449
rect 563501 493374 563513 493408
rect 563547 493374 563559 493408
rect 563501 493340 563559 493374
rect 563501 493306 563513 493340
rect 563547 493306 563559 493340
rect 563501 493272 563559 493306
rect 563501 493238 563513 493272
rect 563547 493238 563559 493272
rect 563501 493204 563559 493238
rect 563501 493170 563513 493204
rect 563547 493170 563559 493204
rect 563501 493136 563559 493170
rect 563501 493102 563513 493136
rect 563547 493102 563559 493136
rect 563501 493068 563559 493102
rect 563501 493034 563513 493068
rect 563547 493034 563559 493068
rect 563501 493000 563559 493034
rect 563501 492966 563513 493000
rect 563547 492966 563559 493000
rect 563501 492932 563559 492966
rect 563501 492898 563513 492932
rect 563547 492898 563559 492932
rect 563501 492864 563559 492898
rect 563501 492830 563513 492864
rect 563547 492830 563559 492864
rect 563501 492796 563559 492830
rect 563501 492762 563513 492796
rect 563547 492762 563559 492796
rect 563501 492728 563559 492762
rect 563501 492694 563513 492728
rect 563547 492694 563559 492728
rect 563501 492660 563559 492694
rect 563501 492626 563513 492660
rect 563547 492626 563559 492660
rect 563501 492592 563559 492626
rect 563501 492558 563513 492592
rect 563547 492558 563559 492592
rect 563501 492524 563559 492558
rect 563501 492490 563513 492524
rect 563547 492490 563559 492524
rect 563501 492449 563559 492490
rect 563759 493408 563817 493449
rect 563759 493374 563771 493408
rect 563805 493374 563817 493408
rect 563759 493340 563817 493374
rect 563759 493306 563771 493340
rect 563805 493306 563817 493340
rect 563759 493272 563817 493306
rect 563759 493238 563771 493272
rect 563805 493238 563817 493272
rect 563759 493204 563817 493238
rect 563759 493170 563771 493204
rect 563805 493170 563817 493204
rect 563759 493136 563817 493170
rect 563759 493102 563771 493136
rect 563805 493102 563817 493136
rect 563759 493068 563817 493102
rect 563759 493034 563771 493068
rect 563805 493034 563817 493068
rect 563759 493000 563817 493034
rect 563759 492966 563771 493000
rect 563805 492966 563817 493000
rect 563759 492932 563817 492966
rect 563759 492898 563771 492932
rect 563805 492898 563817 492932
rect 563759 492864 563817 492898
rect 563759 492830 563771 492864
rect 563805 492830 563817 492864
rect 563759 492796 563817 492830
rect 563759 492762 563771 492796
rect 563805 492762 563817 492796
rect 563759 492728 563817 492762
rect 563759 492694 563771 492728
rect 563805 492694 563817 492728
rect 563759 492660 563817 492694
rect 563759 492626 563771 492660
rect 563805 492626 563817 492660
rect 563759 492592 563817 492626
rect 563759 492558 563771 492592
rect 563805 492558 563817 492592
rect 563759 492524 563817 492558
rect 563759 492490 563771 492524
rect 563805 492490 563817 492524
rect 563759 492449 563817 492490
rect 564017 493408 564075 493449
rect 564017 493374 564029 493408
rect 564063 493374 564075 493408
rect 564017 493340 564075 493374
rect 564017 493306 564029 493340
rect 564063 493306 564075 493340
rect 564017 493272 564075 493306
rect 564017 493238 564029 493272
rect 564063 493238 564075 493272
rect 564017 493204 564075 493238
rect 564017 493170 564029 493204
rect 564063 493170 564075 493204
rect 564017 493136 564075 493170
rect 564017 493102 564029 493136
rect 564063 493102 564075 493136
rect 564017 493068 564075 493102
rect 564017 493034 564029 493068
rect 564063 493034 564075 493068
rect 564017 493000 564075 493034
rect 564017 492966 564029 493000
rect 564063 492966 564075 493000
rect 564017 492932 564075 492966
rect 564017 492898 564029 492932
rect 564063 492898 564075 492932
rect 564017 492864 564075 492898
rect 564017 492830 564029 492864
rect 564063 492830 564075 492864
rect 564017 492796 564075 492830
rect 564017 492762 564029 492796
rect 564063 492762 564075 492796
rect 564017 492728 564075 492762
rect 564017 492694 564029 492728
rect 564063 492694 564075 492728
rect 564017 492660 564075 492694
rect 564017 492626 564029 492660
rect 564063 492626 564075 492660
rect 564017 492592 564075 492626
rect 564017 492558 564029 492592
rect 564063 492558 564075 492592
rect 564017 492524 564075 492558
rect 564017 492490 564029 492524
rect 564063 492490 564075 492524
rect 564017 492449 564075 492490
rect 564275 493408 564333 493449
rect 564275 493374 564287 493408
rect 564321 493374 564333 493408
rect 564275 493340 564333 493374
rect 564275 493306 564287 493340
rect 564321 493306 564333 493340
rect 564275 493272 564333 493306
rect 564275 493238 564287 493272
rect 564321 493238 564333 493272
rect 564275 493204 564333 493238
rect 564275 493170 564287 493204
rect 564321 493170 564333 493204
rect 564275 493136 564333 493170
rect 564275 493102 564287 493136
rect 564321 493102 564333 493136
rect 564275 493068 564333 493102
rect 564275 493034 564287 493068
rect 564321 493034 564333 493068
rect 564275 493000 564333 493034
rect 564275 492966 564287 493000
rect 564321 492966 564333 493000
rect 564275 492932 564333 492966
rect 564275 492898 564287 492932
rect 564321 492898 564333 492932
rect 564275 492864 564333 492898
rect 564275 492830 564287 492864
rect 564321 492830 564333 492864
rect 564275 492796 564333 492830
rect 564275 492762 564287 492796
rect 564321 492762 564333 492796
rect 564275 492728 564333 492762
rect 564275 492694 564287 492728
rect 564321 492694 564333 492728
rect 564275 492660 564333 492694
rect 564275 492626 564287 492660
rect 564321 492626 564333 492660
rect 564275 492592 564333 492626
rect 564275 492558 564287 492592
rect 564321 492558 564333 492592
rect 564275 492524 564333 492558
rect 564275 492490 564287 492524
rect 564321 492490 564333 492524
rect 564275 492449 564333 492490
rect 564533 493408 564591 493449
rect 564533 493374 564545 493408
rect 564579 493374 564591 493408
rect 564533 493340 564591 493374
rect 564533 493306 564545 493340
rect 564579 493306 564591 493340
rect 564533 493272 564591 493306
rect 564533 493238 564545 493272
rect 564579 493238 564591 493272
rect 564533 493204 564591 493238
rect 564533 493170 564545 493204
rect 564579 493170 564591 493204
rect 564533 493136 564591 493170
rect 564533 493102 564545 493136
rect 564579 493102 564591 493136
rect 564533 493068 564591 493102
rect 564533 493034 564545 493068
rect 564579 493034 564591 493068
rect 564533 493000 564591 493034
rect 564533 492966 564545 493000
rect 564579 492966 564591 493000
rect 564533 492932 564591 492966
rect 564533 492898 564545 492932
rect 564579 492898 564591 492932
rect 564533 492864 564591 492898
rect 564533 492830 564545 492864
rect 564579 492830 564591 492864
rect 564533 492796 564591 492830
rect 564533 492762 564545 492796
rect 564579 492762 564591 492796
rect 564533 492728 564591 492762
rect 564533 492694 564545 492728
rect 564579 492694 564591 492728
rect 564533 492660 564591 492694
rect 564533 492626 564545 492660
rect 564579 492626 564591 492660
rect 564533 492592 564591 492626
rect 564533 492558 564545 492592
rect 564579 492558 564591 492592
rect 564533 492524 564591 492558
rect 564533 492490 564545 492524
rect 564579 492490 564591 492524
rect 564533 492449 564591 492490
rect 564791 493408 564849 493449
rect 564791 493374 564803 493408
rect 564837 493374 564849 493408
rect 564791 493340 564849 493374
rect 564791 493306 564803 493340
rect 564837 493306 564849 493340
rect 564791 493272 564849 493306
rect 564791 493238 564803 493272
rect 564837 493238 564849 493272
rect 564791 493204 564849 493238
rect 564791 493170 564803 493204
rect 564837 493170 564849 493204
rect 564791 493136 564849 493170
rect 564791 493102 564803 493136
rect 564837 493102 564849 493136
rect 564791 493068 564849 493102
rect 564791 493034 564803 493068
rect 564837 493034 564849 493068
rect 564791 493000 564849 493034
rect 564791 492966 564803 493000
rect 564837 492966 564849 493000
rect 564791 492932 564849 492966
rect 564791 492898 564803 492932
rect 564837 492898 564849 492932
rect 564791 492864 564849 492898
rect 564791 492830 564803 492864
rect 564837 492830 564849 492864
rect 564791 492796 564849 492830
rect 564791 492762 564803 492796
rect 564837 492762 564849 492796
rect 564791 492728 564849 492762
rect 564791 492694 564803 492728
rect 564837 492694 564849 492728
rect 564791 492660 564849 492694
rect 564791 492626 564803 492660
rect 564837 492626 564849 492660
rect 564791 492592 564849 492626
rect 564791 492558 564803 492592
rect 564837 492558 564849 492592
rect 564791 492524 564849 492558
rect 564791 492490 564803 492524
rect 564837 492490 564849 492524
rect 564791 492449 564849 492490
rect 565049 493408 565107 493449
rect 565049 493374 565061 493408
rect 565095 493374 565107 493408
rect 565049 493340 565107 493374
rect 565049 493306 565061 493340
rect 565095 493306 565107 493340
rect 565049 493272 565107 493306
rect 565049 493238 565061 493272
rect 565095 493238 565107 493272
rect 565049 493204 565107 493238
rect 565049 493170 565061 493204
rect 565095 493170 565107 493204
rect 565049 493136 565107 493170
rect 565049 493102 565061 493136
rect 565095 493102 565107 493136
rect 565049 493068 565107 493102
rect 565049 493034 565061 493068
rect 565095 493034 565107 493068
rect 565049 493000 565107 493034
rect 565049 492966 565061 493000
rect 565095 492966 565107 493000
rect 565049 492932 565107 492966
rect 565049 492898 565061 492932
rect 565095 492898 565107 492932
rect 565049 492864 565107 492898
rect 565049 492830 565061 492864
rect 565095 492830 565107 492864
rect 565049 492796 565107 492830
rect 565049 492762 565061 492796
rect 565095 492762 565107 492796
rect 565049 492728 565107 492762
rect 565049 492694 565061 492728
rect 565095 492694 565107 492728
rect 565049 492660 565107 492694
rect 565049 492626 565061 492660
rect 565095 492626 565107 492660
rect 565049 492592 565107 492626
rect 565049 492558 565061 492592
rect 565095 492558 565107 492592
rect 565049 492524 565107 492558
rect 565049 492490 565061 492524
rect 565095 492490 565107 492524
rect 565049 492449 565107 492490
rect 565307 493408 565365 493449
rect 565307 493374 565319 493408
rect 565353 493374 565365 493408
rect 565307 493340 565365 493374
rect 565307 493306 565319 493340
rect 565353 493306 565365 493340
rect 565307 493272 565365 493306
rect 565307 493238 565319 493272
rect 565353 493238 565365 493272
rect 565307 493204 565365 493238
rect 565307 493170 565319 493204
rect 565353 493170 565365 493204
rect 565307 493136 565365 493170
rect 565307 493102 565319 493136
rect 565353 493102 565365 493136
rect 565307 493068 565365 493102
rect 565307 493034 565319 493068
rect 565353 493034 565365 493068
rect 565307 493000 565365 493034
rect 565307 492966 565319 493000
rect 565353 492966 565365 493000
rect 565307 492932 565365 492966
rect 565307 492898 565319 492932
rect 565353 492898 565365 492932
rect 565307 492864 565365 492898
rect 565307 492830 565319 492864
rect 565353 492830 565365 492864
rect 565307 492796 565365 492830
rect 565307 492762 565319 492796
rect 565353 492762 565365 492796
rect 565307 492728 565365 492762
rect 565307 492694 565319 492728
rect 565353 492694 565365 492728
rect 565307 492660 565365 492694
rect 565307 492626 565319 492660
rect 565353 492626 565365 492660
rect 565307 492592 565365 492626
rect 565307 492558 565319 492592
rect 565353 492558 565365 492592
rect 565307 492524 565365 492558
rect 565307 492490 565319 492524
rect 565353 492490 565365 492524
rect 565307 492449 565365 492490
rect 565565 493408 565623 493449
rect 565565 493374 565577 493408
rect 565611 493374 565623 493408
rect 565565 493340 565623 493374
rect 565565 493306 565577 493340
rect 565611 493306 565623 493340
rect 565565 493272 565623 493306
rect 565565 493238 565577 493272
rect 565611 493238 565623 493272
rect 565565 493204 565623 493238
rect 565565 493170 565577 493204
rect 565611 493170 565623 493204
rect 565565 493136 565623 493170
rect 565565 493102 565577 493136
rect 565611 493102 565623 493136
rect 565565 493068 565623 493102
rect 565565 493034 565577 493068
rect 565611 493034 565623 493068
rect 565565 493000 565623 493034
rect 565565 492966 565577 493000
rect 565611 492966 565623 493000
rect 565565 492932 565623 492966
rect 565565 492898 565577 492932
rect 565611 492898 565623 492932
rect 565565 492864 565623 492898
rect 565565 492830 565577 492864
rect 565611 492830 565623 492864
rect 565565 492796 565623 492830
rect 565565 492762 565577 492796
rect 565611 492762 565623 492796
rect 565565 492728 565623 492762
rect 565565 492694 565577 492728
rect 565611 492694 565623 492728
rect 565565 492660 565623 492694
rect 565565 492626 565577 492660
rect 565611 492626 565623 492660
rect 565565 492592 565623 492626
rect 565565 492558 565577 492592
rect 565611 492558 565623 492592
rect 565565 492524 565623 492558
rect 565565 492490 565577 492524
rect 565611 492490 565623 492524
rect 565565 492449 565623 492490
rect 565823 493408 565881 493449
rect 565823 493374 565835 493408
rect 565869 493374 565881 493408
rect 565823 493340 565881 493374
rect 565823 493306 565835 493340
rect 565869 493306 565881 493340
rect 565823 493272 565881 493306
rect 565823 493238 565835 493272
rect 565869 493238 565881 493272
rect 565823 493204 565881 493238
rect 565823 493170 565835 493204
rect 565869 493170 565881 493204
rect 565823 493136 565881 493170
rect 565823 493102 565835 493136
rect 565869 493102 565881 493136
rect 565823 493068 565881 493102
rect 565823 493034 565835 493068
rect 565869 493034 565881 493068
rect 565823 493000 565881 493034
rect 565823 492966 565835 493000
rect 565869 492966 565881 493000
rect 565823 492932 565881 492966
rect 565823 492898 565835 492932
rect 565869 492898 565881 492932
rect 565823 492864 565881 492898
rect 565823 492830 565835 492864
rect 565869 492830 565881 492864
rect 565823 492796 565881 492830
rect 565823 492762 565835 492796
rect 565869 492762 565881 492796
rect 565823 492728 565881 492762
rect 565823 492694 565835 492728
rect 565869 492694 565881 492728
rect 565823 492660 565881 492694
rect 565823 492626 565835 492660
rect 565869 492626 565881 492660
rect 565823 492592 565881 492626
rect 565823 492558 565835 492592
rect 565869 492558 565881 492592
rect 565823 492524 565881 492558
rect 565823 492490 565835 492524
rect 565869 492490 565881 492524
rect 565823 492449 565881 492490
rect 560599 404266 560657 404307
rect 560599 404232 560611 404266
rect 560645 404232 560657 404266
rect 560599 404198 560657 404232
rect 560599 404164 560611 404198
rect 560645 404164 560657 404198
rect 560599 404130 560657 404164
rect 560599 404096 560611 404130
rect 560645 404096 560657 404130
rect 560599 404062 560657 404096
rect 560599 404028 560611 404062
rect 560645 404028 560657 404062
rect 560599 403994 560657 404028
rect 560599 403960 560611 403994
rect 560645 403960 560657 403994
rect 560599 403926 560657 403960
rect 560599 403892 560611 403926
rect 560645 403892 560657 403926
rect 560599 403858 560657 403892
rect 560599 403824 560611 403858
rect 560645 403824 560657 403858
rect 560599 403790 560657 403824
rect 560599 403756 560611 403790
rect 560645 403756 560657 403790
rect 560599 403722 560657 403756
rect 560599 403688 560611 403722
rect 560645 403688 560657 403722
rect 560599 403654 560657 403688
rect 560599 403620 560611 403654
rect 560645 403620 560657 403654
rect 560599 403586 560657 403620
rect 560599 403552 560611 403586
rect 560645 403552 560657 403586
rect 560599 403518 560657 403552
rect 560599 403484 560611 403518
rect 560645 403484 560657 403518
rect 560599 403450 560657 403484
rect 560599 403416 560611 403450
rect 560645 403416 560657 403450
rect 560599 403382 560657 403416
rect 560599 403348 560611 403382
rect 560645 403348 560657 403382
rect 560599 403307 560657 403348
rect 560857 404266 560915 404307
rect 560857 404232 560869 404266
rect 560903 404232 560915 404266
rect 560857 404198 560915 404232
rect 560857 404164 560869 404198
rect 560903 404164 560915 404198
rect 560857 404130 560915 404164
rect 560857 404096 560869 404130
rect 560903 404096 560915 404130
rect 560857 404062 560915 404096
rect 560857 404028 560869 404062
rect 560903 404028 560915 404062
rect 560857 403994 560915 404028
rect 560857 403960 560869 403994
rect 560903 403960 560915 403994
rect 560857 403926 560915 403960
rect 560857 403892 560869 403926
rect 560903 403892 560915 403926
rect 560857 403858 560915 403892
rect 560857 403824 560869 403858
rect 560903 403824 560915 403858
rect 560857 403790 560915 403824
rect 560857 403756 560869 403790
rect 560903 403756 560915 403790
rect 560857 403722 560915 403756
rect 560857 403688 560869 403722
rect 560903 403688 560915 403722
rect 560857 403654 560915 403688
rect 560857 403620 560869 403654
rect 560903 403620 560915 403654
rect 560857 403586 560915 403620
rect 560857 403552 560869 403586
rect 560903 403552 560915 403586
rect 560857 403518 560915 403552
rect 560857 403484 560869 403518
rect 560903 403484 560915 403518
rect 560857 403450 560915 403484
rect 560857 403416 560869 403450
rect 560903 403416 560915 403450
rect 560857 403382 560915 403416
rect 560857 403348 560869 403382
rect 560903 403348 560915 403382
rect 560857 403307 560915 403348
rect 561115 404266 561173 404307
rect 561115 404232 561127 404266
rect 561161 404232 561173 404266
rect 561115 404198 561173 404232
rect 561115 404164 561127 404198
rect 561161 404164 561173 404198
rect 561115 404130 561173 404164
rect 561115 404096 561127 404130
rect 561161 404096 561173 404130
rect 561115 404062 561173 404096
rect 561115 404028 561127 404062
rect 561161 404028 561173 404062
rect 561115 403994 561173 404028
rect 561115 403960 561127 403994
rect 561161 403960 561173 403994
rect 561115 403926 561173 403960
rect 561115 403892 561127 403926
rect 561161 403892 561173 403926
rect 561115 403858 561173 403892
rect 561115 403824 561127 403858
rect 561161 403824 561173 403858
rect 561115 403790 561173 403824
rect 561115 403756 561127 403790
rect 561161 403756 561173 403790
rect 561115 403722 561173 403756
rect 561115 403688 561127 403722
rect 561161 403688 561173 403722
rect 561115 403654 561173 403688
rect 561115 403620 561127 403654
rect 561161 403620 561173 403654
rect 561115 403586 561173 403620
rect 561115 403552 561127 403586
rect 561161 403552 561173 403586
rect 561115 403518 561173 403552
rect 561115 403484 561127 403518
rect 561161 403484 561173 403518
rect 561115 403450 561173 403484
rect 561115 403416 561127 403450
rect 561161 403416 561173 403450
rect 561115 403382 561173 403416
rect 561115 403348 561127 403382
rect 561161 403348 561173 403382
rect 561115 403307 561173 403348
rect 561373 404266 561431 404307
rect 561373 404232 561385 404266
rect 561419 404232 561431 404266
rect 561373 404198 561431 404232
rect 561373 404164 561385 404198
rect 561419 404164 561431 404198
rect 561373 404130 561431 404164
rect 561373 404096 561385 404130
rect 561419 404096 561431 404130
rect 561373 404062 561431 404096
rect 561373 404028 561385 404062
rect 561419 404028 561431 404062
rect 561373 403994 561431 404028
rect 561373 403960 561385 403994
rect 561419 403960 561431 403994
rect 561373 403926 561431 403960
rect 561373 403892 561385 403926
rect 561419 403892 561431 403926
rect 561373 403858 561431 403892
rect 561373 403824 561385 403858
rect 561419 403824 561431 403858
rect 561373 403790 561431 403824
rect 561373 403756 561385 403790
rect 561419 403756 561431 403790
rect 561373 403722 561431 403756
rect 561373 403688 561385 403722
rect 561419 403688 561431 403722
rect 561373 403654 561431 403688
rect 561373 403620 561385 403654
rect 561419 403620 561431 403654
rect 561373 403586 561431 403620
rect 561373 403552 561385 403586
rect 561419 403552 561431 403586
rect 561373 403518 561431 403552
rect 561373 403484 561385 403518
rect 561419 403484 561431 403518
rect 561373 403450 561431 403484
rect 561373 403416 561385 403450
rect 561419 403416 561431 403450
rect 561373 403382 561431 403416
rect 561373 403348 561385 403382
rect 561419 403348 561431 403382
rect 561373 403307 561431 403348
rect 561631 404266 561689 404307
rect 561631 404232 561643 404266
rect 561677 404232 561689 404266
rect 561631 404198 561689 404232
rect 561631 404164 561643 404198
rect 561677 404164 561689 404198
rect 561631 404130 561689 404164
rect 561631 404096 561643 404130
rect 561677 404096 561689 404130
rect 561631 404062 561689 404096
rect 561631 404028 561643 404062
rect 561677 404028 561689 404062
rect 561631 403994 561689 404028
rect 561631 403960 561643 403994
rect 561677 403960 561689 403994
rect 561631 403926 561689 403960
rect 561631 403892 561643 403926
rect 561677 403892 561689 403926
rect 561631 403858 561689 403892
rect 561631 403824 561643 403858
rect 561677 403824 561689 403858
rect 561631 403790 561689 403824
rect 561631 403756 561643 403790
rect 561677 403756 561689 403790
rect 561631 403722 561689 403756
rect 561631 403688 561643 403722
rect 561677 403688 561689 403722
rect 561631 403654 561689 403688
rect 561631 403620 561643 403654
rect 561677 403620 561689 403654
rect 561631 403586 561689 403620
rect 561631 403552 561643 403586
rect 561677 403552 561689 403586
rect 561631 403518 561689 403552
rect 561631 403484 561643 403518
rect 561677 403484 561689 403518
rect 561631 403450 561689 403484
rect 561631 403416 561643 403450
rect 561677 403416 561689 403450
rect 561631 403382 561689 403416
rect 561631 403348 561643 403382
rect 561677 403348 561689 403382
rect 561631 403307 561689 403348
rect 561889 404266 561947 404307
rect 561889 404232 561901 404266
rect 561935 404232 561947 404266
rect 561889 404198 561947 404232
rect 561889 404164 561901 404198
rect 561935 404164 561947 404198
rect 561889 404130 561947 404164
rect 561889 404096 561901 404130
rect 561935 404096 561947 404130
rect 561889 404062 561947 404096
rect 561889 404028 561901 404062
rect 561935 404028 561947 404062
rect 561889 403994 561947 404028
rect 561889 403960 561901 403994
rect 561935 403960 561947 403994
rect 561889 403926 561947 403960
rect 561889 403892 561901 403926
rect 561935 403892 561947 403926
rect 561889 403858 561947 403892
rect 561889 403824 561901 403858
rect 561935 403824 561947 403858
rect 561889 403790 561947 403824
rect 561889 403756 561901 403790
rect 561935 403756 561947 403790
rect 561889 403722 561947 403756
rect 561889 403688 561901 403722
rect 561935 403688 561947 403722
rect 561889 403654 561947 403688
rect 561889 403620 561901 403654
rect 561935 403620 561947 403654
rect 561889 403586 561947 403620
rect 561889 403552 561901 403586
rect 561935 403552 561947 403586
rect 561889 403518 561947 403552
rect 561889 403484 561901 403518
rect 561935 403484 561947 403518
rect 561889 403450 561947 403484
rect 561889 403416 561901 403450
rect 561935 403416 561947 403450
rect 561889 403382 561947 403416
rect 561889 403348 561901 403382
rect 561935 403348 561947 403382
rect 561889 403307 561947 403348
rect 562147 404266 562205 404307
rect 562147 404232 562159 404266
rect 562193 404232 562205 404266
rect 562147 404198 562205 404232
rect 562147 404164 562159 404198
rect 562193 404164 562205 404198
rect 562147 404130 562205 404164
rect 562147 404096 562159 404130
rect 562193 404096 562205 404130
rect 562147 404062 562205 404096
rect 562147 404028 562159 404062
rect 562193 404028 562205 404062
rect 562147 403994 562205 404028
rect 562147 403960 562159 403994
rect 562193 403960 562205 403994
rect 562147 403926 562205 403960
rect 562147 403892 562159 403926
rect 562193 403892 562205 403926
rect 562147 403858 562205 403892
rect 562147 403824 562159 403858
rect 562193 403824 562205 403858
rect 562147 403790 562205 403824
rect 562147 403756 562159 403790
rect 562193 403756 562205 403790
rect 562147 403722 562205 403756
rect 562147 403688 562159 403722
rect 562193 403688 562205 403722
rect 562147 403654 562205 403688
rect 562147 403620 562159 403654
rect 562193 403620 562205 403654
rect 562147 403586 562205 403620
rect 562147 403552 562159 403586
rect 562193 403552 562205 403586
rect 562147 403518 562205 403552
rect 562147 403484 562159 403518
rect 562193 403484 562205 403518
rect 562147 403450 562205 403484
rect 562147 403416 562159 403450
rect 562193 403416 562205 403450
rect 562147 403382 562205 403416
rect 562147 403348 562159 403382
rect 562193 403348 562205 403382
rect 562147 403307 562205 403348
rect 562405 404266 562463 404307
rect 562405 404232 562417 404266
rect 562451 404232 562463 404266
rect 562405 404198 562463 404232
rect 562405 404164 562417 404198
rect 562451 404164 562463 404198
rect 562405 404130 562463 404164
rect 562405 404096 562417 404130
rect 562451 404096 562463 404130
rect 562405 404062 562463 404096
rect 562405 404028 562417 404062
rect 562451 404028 562463 404062
rect 562405 403994 562463 404028
rect 562405 403960 562417 403994
rect 562451 403960 562463 403994
rect 562405 403926 562463 403960
rect 562405 403892 562417 403926
rect 562451 403892 562463 403926
rect 562405 403858 562463 403892
rect 562405 403824 562417 403858
rect 562451 403824 562463 403858
rect 562405 403790 562463 403824
rect 562405 403756 562417 403790
rect 562451 403756 562463 403790
rect 562405 403722 562463 403756
rect 562405 403688 562417 403722
rect 562451 403688 562463 403722
rect 562405 403654 562463 403688
rect 562405 403620 562417 403654
rect 562451 403620 562463 403654
rect 562405 403586 562463 403620
rect 562405 403552 562417 403586
rect 562451 403552 562463 403586
rect 562405 403518 562463 403552
rect 562405 403484 562417 403518
rect 562451 403484 562463 403518
rect 562405 403450 562463 403484
rect 562405 403416 562417 403450
rect 562451 403416 562463 403450
rect 562405 403382 562463 403416
rect 562405 403348 562417 403382
rect 562451 403348 562463 403382
rect 562405 403307 562463 403348
rect 562663 404266 562721 404307
rect 562663 404232 562675 404266
rect 562709 404232 562721 404266
rect 562663 404198 562721 404232
rect 562663 404164 562675 404198
rect 562709 404164 562721 404198
rect 562663 404130 562721 404164
rect 562663 404096 562675 404130
rect 562709 404096 562721 404130
rect 562663 404062 562721 404096
rect 562663 404028 562675 404062
rect 562709 404028 562721 404062
rect 562663 403994 562721 404028
rect 562663 403960 562675 403994
rect 562709 403960 562721 403994
rect 562663 403926 562721 403960
rect 562663 403892 562675 403926
rect 562709 403892 562721 403926
rect 562663 403858 562721 403892
rect 562663 403824 562675 403858
rect 562709 403824 562721 403858
rect 562663 403790 562721 403824
rect 562663 403756 562675 403790
rect 562709 403756 562721 403790
rect 562663 403722 562721 403756
rect 562663 403688 562675 403722
rect 562709 403688 562721 403722
rect 562663 403654 562721 403688
rect 562663 403620 562675 403654
rect 562709 403620 562721 403654
rect 562663 403586 562721 403620
rect 562663 403552 562675 403586
rect 562709 403552 562721 403586
rect 562663 403518 562721 403552
rect 562663 403484 562675 403518
rect 562709 403484 562721 403518
rect 562663 403450 562721 403484
rect 562663 403416 562675 403450
rect 562709 403416 562721 403450
rect 562663 403382 562721 403416
rect 562663 403348 562675 403382
rect 562709 403348 562721 403382
rect 562663 403307 562721 403348
rect 562921 404266 562979 404307
rect 562921 404232 562933 404266
rect 562967 404232 562979 404266
rect 562921 404198 562979 404232
rect 562921 404164 562933 404198
rect 562967 404164 562979 404198
rect 562921 404130 562979 404164
rect 562921 404096 562933 404130
rect 562967 404096 562979 404130
rect 562921 404062 562979 404096
rect 562921 404028 562933 404062
rect 562967 404028 562979 404062
rect 562921 403994 562979 404028
rect 562921 403960 562933 403994
rect 562967 403960 562979 403994
rect 562921 403926 562979 403960
rect 562921 403892 562933 403926
rect 562967 403892 562979 403926
rect 562921 403858 562979 403892
rect 562921 403824 562933 403858
rect 562967 403824 562979 403858
rect 562921 403790 562979 403824
rect 562921 403756 562933 403790
rect 562967 403756 562979 403790
rect 562921 403722 562979 403756
rect 562921 403688 562933 403722
rect 562967 403688 562979 403722
rect 562921 403654 562979 403688
rect 562921 403620 562933 403654
rect 562967 403620 562979 403654
rect 562921 403586 562979 403620
rect 562921 403552 562933 403586
rect 562967 403552 562979 403586
rect 562921 403518 562979 403552
rect 562921 403484 562933 403518
rect 562967 403484 562979 403518
rect 562921 403450 562979 403484
rect 562921 403416 562933 403450
rect 562967 403416 562979 403450
rect 562921 403382 562979 403416
rect 562921 403348 562933 403382
rect 562967 403348 562979 403382
rect 562921 403307 562979 403348
rect 563179 404266 563237 404307
rect 563179 404232 563191 404266
rect 563225 404232 563237 404266
rect 563179 404198 563237 404232
rect 563179 404164 563191 404198
rect 563225 404164 563237 404198
rect 563179 404130 563237 404164
rect 563179 404096 563191 404130
rect 563225 404096 563237 404130
rect 563179 404062 563237 404096
rect 563179 404028 563191 404062
rect 563225 404028 563237 404062
rect 563179 403994 563237 404028
rect 563179 403960 563191 403994
rect 563225 403960 563237 403994
rect 563179 403926 563237 403960
rect 563179 403892 563191 403926
rect 563225 403892 563237 403926
rect 563179 403858 563237 403892
rect 563179 403824 563191 403858
rect 563225 403824 563237 403858
rect 563179 403790 563237 403824
rect 563179 403756 563191 403790
rect 563225 403756 563237 403790
rect 563179 403722 563237 403756
rect 563179 403688 563191 403722
rect 563225 403688 563237 403722
rect 563179 403654 563237 403688
rect 563179 403620 563191 403654
rect 563225 403620 563237 403654
rect 563179 403586 563237 403620
rect 563179 403552 563191 403586
rect 563225 403552 563237 403586
rect 563179 403518 563237 403552
rect 563179 403484 563191 403518
rect 563225 403484 563237 403518
rect 563179 403450 563237 403484
rect 563179 403416 563191 403450
rect 563225 403416 563237 403450
rect 563179 403382 563237 403416
rect 563179 403348 563191 403382
rect 563225 403348 563237 403382
rect 563179 403307 563237 403348
rect 563437 404266 563495 404307
rect 563437 404232 563449 404266
rect 563483 404232 563495 404266
rect 563437 404198 563495 404232
rect 563437 404164 563449 404198
rect 563483 404164 563495 404198
rect 563437 404130 563495 404164
rect 563437 404096 563449 404130
rect 563483 404096 563495 404130
rect 563437 404062 563495 404096
rect 563437 404028 563449 404062
rect 563483 404028 563495 404062
rect 563437 403994 563495 404028
rect 563437 403960 563449 403994
rect 563483 403960 563495 403994
rect 563437 403926 563495 403960
rect 563437 403892 563449 403926
rect 563483 403892 563495 403926
rect 563437 403858 563495 403892
rect 563437 403824 563449 403858
rect 563483 403824 563495 403858
rect 563437 403790 563495 403824
rect 563437 403756 563449 403790
rect 563483 403756 563495 403790
rect 563437 403722 563495 403756
rect 563437 403688 563449 403722
rect 563483 403688 563495 403722
rect 563437 403654 563495 403688
rect 563437 403620 563449 403654
rect 563483 403620 563495 403654
rect 563437 403586 563495 403620
rect 563437 403552 563449 403586
rect 563483 403552 563495 403586
rect 563437 403518 563495 403552
rect 563437 403484 563449 403518
rect 563483 403484 563495 403518
rect 563437 403450 563495 403484
rect 563437 403416 563449 403450
rect 563483 403416 563495 403450
rect 563437 403382 563495 403416
rect 563437 403348 563449 403382
rect 563483 403348 563495 403382
rect 563437 403307 563495 403348
rect 563695 404266 563753 404307
rect 563695 404232 563707 404266
rect 563741 404232 563753 404266
rect 563695 404198 563753 404232
rect 563695 404164 563707 404198
rect 563741 404164 563753 404198
rect 563695 404130 563753 404164
rect 563695 404096 563707 404130
rect 563741 404096 563753 404130
rect 563695 404062 563753 404096
rect 563695 404028 563707 404062
rect 563741 404028 563753 404062
rect 563695 403994 563753 404028
rect 563695 403960 563707 403994
rect 563741 403960 563753 403994
rect 563695 403926 563753 403960
rect 563695 403892 563707 403926
rect 563741 403892 563753 403926
rect 563695 403858 563753 403892
rect 563695 403824 563707 403858
rect 563741 403824 563753 403858
rect 563695 403790 563753 403824
rect 563695 403756 563707 403790
rect 563741 403756 563753 403790
rect 563695 403722 563753 403756
rect 563695 403688 563707 403722
rect 563741 403688 563753 403722
rect 563695 403654 563753 403688
rect 563695 403620 563707 403654
rect 563741 403620 563753 403654
rect 563695 403586 563753 403620
rect 563695 403552 563707 403586
rect 563741 403552 563753 403586
rect 563695 403518 563753 403552
rect 563695 403484 563707 403518
rect 563741 403484 563753 403518
rect 563695 403450 563753 403484
rect 563695 403416 563707 403450
rect 563741 403416 563753 403450
rect 563695 403382 563753 403416
rect 563695 403348 563707 403382
rect 563741 403348 563753 403382
rect 563695 403307 563753 403348
rect 563953 404266 564011 404307
rect 563953 404232 563965 404266
rect 563999 404232 564011 404266
rect 563953 404198 564011 404232
rect 563953 404164 563965 404198
rect 563999 404164 564011 404198
rect 563953 404130 564011 404164
rect 563953 404096 563965 404130
rect 563999 404096 564011 404130
rect 563953 404062 564011 404096
rect 563953 404028 563965 404062
rect 563999 404028 564011 404062
rect 563953 403994 564011 404028
rect 563953 403960 563965 403994
rect 563999 403960 564011 403994
rect 563953 403926 564011 403960
rect 563953 403892 563965 403926
rect 563999 403892 564011 403926
rect 563953 403858 564011 403892
rect 563953 403824 563965 403858
rect 563999 403824 564011 403858
rect 563953 403790 564011 403824
rect 563953 403756 563965 403790
rect 563999 403756 564011 403790
rect 563953 403722 564011 403756
rect 563953 403688 563965 403722
rect 563999 403688 564011 403722
rect 563953 403654 564011 403688
rect 563953 403620 563965 403654
rect 563999 403620 564011 403654
rect 563953 403586 564011 403620
rect 563953 403552 563965 403586
rect 563999 403552 564011 403586
rect 563953 403518 564011 403552
rect 563953 403484 563965 403518
rect 563999 403484 564011 403518
rect 563953 403450 564011 403484
rect 563953 403416 563965 403450
rect 563999 403416 564011 403450
rect 563953 403382 564011 403416
rect 563953 403348 563965 403382
rect 563999 403348 564011 403382
rect 563953 403307 564011 403348
rect 564211 404266 564269 404307
rect 564211 404232 564223 404266
rect 564257 404232 564269 404266
rect 564211 404198 564269 404232
rect 564211 404164 564223 404198
rect 564257 404164 564269 404198
rect 564211 404130 564269 404164
rect 564211 404096 564223 404130
rect 564257 404096 564269 404130
rect 564211 404062 564269 404096
rect 564211 404028 564223 404062
rect 564257 404028 564269 404062
rect 564211 403994 564269 404028
rect 564211 403960 564223 403994
rect 564257 403960 564269 403994
rect 564211 403926 564269 403960
rect 564211 403892 564223 403926
rect 564257 403892 564269 403926
rect 564211 403858 564269 403892
rect 564211 403824 564223 403858
rect 564257 403824 564269 403858
rect 564211 403790 564269 403824
rect 564211 403756 564223 403790
rect 564257 403756 564269 403790
rect 564211 403722 564269 403756
rect 564211 403688 564223 403722
rect 564257 403688 564269 403722
rect 564211 403654 564269 403688
rect 564211 403620 564223 403654
rect 564257 403620 564269 403654
rect 564211 403586 564269 403620
rect 564211 403552 564223 403586
rect 564257 403552 564269 403586
rect 564211 403518 564269 403552
rect 564211 403484 564223 403518
rect 564257 403484 564269 403518
rect 564211 403450 564269 403484
rect 564211 403416 564223 403450
rect 564257 403416 564269 403450
rect 564211 403382 564269 403416
rect 564211 403348 564223 403382
rect 564257 403348 564269 403382
rect 564211 403307 564269 403348
rect 564469 404266 564527 404307
rect 564469 404232 564481 404266
rect 564515 404232 564527 404266
rect 564469 404198 564527 404232
rect 564469 404164 564481 404198
rect 564515 404164 564527 404198
rect 564469 404130 564527 404164
rect 564469 404096 564481 404130
rect 564515 404096 564527 404130
rect 564469 404062 564527 404096
rect 564469 404028 564481 404062
rect 564515 404028 564527 404062
rect 564469 403994 564527 404028
rect 564469 403960 564481 403994
rect 564515 403960 564527 403994
rect 564469 403926 564527 403960
rect 564469 403892 564481 403926
rect 564515 403892 564527 403926
rect 564469 403858 564527 403892
rect 564469 403824 564481 403858
rect 564515 403824 564527 403858
rect 564469 403790 564527 403824
rect 564469 403756 564481 403790
rect 564515 403756 564527 403790
rect 564469 403722 564527 403756
rect 564469 403688 564481 403722
rect 564515 403688 564527 403722
rect 564469 403654 564527 403688
rect 564469 403620 564481 403654
rect 564515 403620 564527 403654
rect 564469 403586 564527 403620
rect 564469 403552 564481 403586
rect 564515 403552 564527 403586
rect 564469 403518 564527 403552
rect 564469 403484 564481 403518
rect 564515 403484 564527 403518
rect 564469 403450 564527 403484
rect 564469 403416 564481 403450
rect 564515 403416 564527 403450
rect 564469 403382 564527 403416
rect 564469 403348 564481 403382
rect 564515 403348 564527 403382
rect 564469 403307 564527 403348
rect 564727 404266 564785 404307
rect 564727 404232 564739 404266
rect 564773 404232 564785 404266
rect 564727 404198 564785 404232
rect 564727 404164 564739 404198
rect 564773 404164 564785 404198
rect 564727 404130 564785 404164
rect 564727 404096 564739 404130
rect 564773 404096 564785 404130
rect 564727 404062 564785 404096
rect 564727 404028 564739 404062
rect 564773 404028 564785 404062
rect 564727 403994 564785 404028
rect 564727 403960 564739 403994
rect 564773 403960 564785 403994
rect 564727 403926 564785 403960
rect 564727 403892 564739 403926
rect 564773 403892 564785 403926
rect 564727 403858 564785 403892
rect 564727 403824 564739 403858
rect 564773 403824 564785 403858
rect 564727 403790 564785 403824
rect 564727 403756 564739 403790
rect 564773 403756 564785 403790
rect 564727 403722 564785 403756
rect 564727 403688 564739 403722
rect 564773 403688 564785 403722
rect 564727 403654 564785 403688
rect 564727 403620 564739 403654
rect 564773 403620 564785 403654
rect 564727 403586 564785 403620
rect 564727 403552 564739 403586
rect 564773 403552 564785 403586
rect 564727 403518 564785 403552
rect 564727 403484 564739 403518
rect 564773 403484 564785 403518
rect 564727 403450 564785 403484
rect 564727 403416 564739 403450
rect 564773 403416 564785 403450
rect 564727 403382 564785 403416
rect 564727 403348 564739 403382
rect 564773 403348 564785 403382
rect 564727 403307 564785 403348
rect 564985 404266 565043 404307
rect 564985 404232 564997 404266
rect 565031 404232 565043 404266
rect 564985 404198 565043 404232
rect 564985 404164 564997 404198
rect 565031 404164 565043 404198
rect 564985 404130 565043 404164
rect 564985 404096 564997 404130
rect 565031 404096 565043 404130
rect 564985 404062 565043 404096
rect 564985 404028 564997 404062
rect 565031 404028 565043 404062
rect 564985 403994 565043 404028
rect 564985 403960 564997 403994
rect 565031 403960 565043 403994
rect 564985 403926 565043 403960
rect 564985 403892 564997 403926
rect 565031 403892 565043 403926
rect 564985 403858 565043 403892
rect 564985 403824 564997 403858
rect 565031 403824 565043 403858
rect 564985 403790 565043 403824
rect 564985 403756 564997 403790
rect 565031 403756 565043 403790
rect 564985 403722 565043 403756
rect 564985 403688 564997 403722
rect 565031 403688 565043 403722
rect 564985 403654 565043 403688
rect 564985 403620 564997 403654
rect 565031 403620 565043 403654
rect 564985 403586 565043 403620
rect 564985 403552 564997 403586
rect 565031 403552 565043 403586
rect 564985 403518 565043 403552
rect 564985 403484 564997 403518
rect 565031 403484 565043 403518
rect 564985 403450 565043 403484
rect 564985 403416 564997 403450
rect 565031 403416 565043 403450
rect 564985 403382 565043 403416
rect 564985 403348 564997 403382
rect 565031 403348 565043 403382
rect 564985 403307 565043 403348
rect 565243 404266 565301 404307
rect 565243 404232 565255 404266
rect 565289 404232 565301 404266
rect 565243 404198 565301 404232
rect 565243 404164 565255 404198
rect 565289 404164 565301 404198
rect 565243 404130 565301 404164
rect 565243 404096 565255 404130
rect 565289 404096 565301 404130
rect 565243 404062 565301 404096
rect 565243 404028 565255 404062
rect 565289 404028 565301 404062
rect 565243 403994 565301 404028
rect 565243 403960 565255 403994
rect 565289 403960 565301 403994
rect 565243 403926 565301 403960
rect 565243 403892 565255 403926
rect 565289 403892 565301 403926
rect 565243 403858 565301 403892
rect 565243 403824 565255 403858
rect 565289 403824 565301 403858
rect 565243 403790 565301 403824
rect 565243 403756 565255 403790
rect 565289 403756 565301 403790
rect 565243 403722 565301 403756
rect 565243 403688 565255 403722
rect 565289 403688 565301 403722
rect 565243 403654 565301 403688
rect 565243 403620 565255 403654
rect 565289 403620 565301 403654
rect 565243 403586 565301 403620
rect 565243 403552 565255 403586
rect 565289 403552 565301 403586
rect 565243 403518 565301 403552
rect 565243 403484 565255 403518
rect 565289 403484 565301 403518
rect 565243 403450 565301 403484
rect 565243 403416 565255 403450
rect 565289 403416 565301 403450
rect 565243 403382 565301 403416
rect 565243 403348 565255 403382
rect 565289 403348 565301 403382
rect 565243 403307 565301 403348
rect 565501 404266 565559 404307
rect 565501 404232 565513 404266
rect 565547 404232 565559 404266
rect 565501 404198 565559 404232
rect 565501 404164 565513 404198
rect 565547 404164 565559 404198
rect 565501 404130 565559 404164
rect 565501 404096 565513 404130
rect 565547 404096 565559 404130
rect 565501 404062 565559 404096
rect 565501 404028 565513 404062
rect 565547 404028 565559 404062
rect 565501 403994 565559 404028
rect 565501 403960 565513 403994
rect 565547 403960 565559 403994
rect 565501 403926 565559 403960
rect 565501 403892 565513 403926
rect 565547 403892 565559 403926
rect 565501 403858 565559 403892
rect 565501 403824 565513 403858
rect 565547 403824 565559 403858
rect 565501 403790 565559 403824
rect 565501 403756 565513 403790
rect 565547 403756 565559 403790
rect 565501 403722 565559 403756
rect 565501 403688 565513 403722
rect 565547 403688 565559 403722
rect 565501 403654 565559 403688
rect 565501 403620 565513 403654
rect 565547 403620 565559 403654
rect 565501 403586 565559 403620
rect 565501 403552 565513 403586
rect 565547 403552 565559 403586
rect 565501 403518 565559 403552
rect 565501 403484 565513 403518
rect 565547 403484 565559 403518
rect 565501 403450 565559 403484
rect 565501 403416 565513 403450
rect 565547 403416 565559 403450
rect 565501 403382 565559 403416
rect 565501 403348 565513 403382
rect 565547 403348 565559 403382
rect 565501 403307 565559 403348
rect 565759 404266 565817 404307
rect 565759 404232 565771 404266
rect 565805 404232 565817 404266
rect 565759 404198 565817 404232
rect 565759 404164 565771 404198
rect 565805 404164 565817 404198
rect 565759 404130 565817 404164
rect 565759 404096 565771 404130
rect 565805 404096 565817 404130
rect 565759 404062 565817 404096
rect 565759 404028 565771 404062
rect 565805 404028 565817 404062
rect 565759 403994 565817 404028
rect 565759 403960 565771 403994
rect 565805 403960 565817 403994
rect 565759 403926 565817 403960
rect 565759 403892 565771 403926
rect 565805 403892 565817 403926
rect 565759 403858 565817 403892
rect 565759 403824 565771 403858
rect 565805 403824 565817 403858
rect 565759 403790 565817 403824
rect 565759 403756 565771 403790
rect 565805 403756 565817 403790
rect 565759 403722 565817 403756
rect 565759 403688 565771 403722
rect 565805 403688 565817 403722
rect 565759 403654 565817 403688
rect 565759 403620 565771 403654
rect 565805 403620 565817 403654
rect 565759 403586 565817 403620
rect 565759 403552 565771 403586
rect 565805 403552 565817 403586
rect 565759 403518 565817 403552
rect 565759 403484 565771 403518
rect 565805 403484 565817 403518
rect 565759 403450 565817 403484
rect 565759 403416 565771 403450
rect 565805 403416 565817 403450
rect 565759 403382 565817 403416
rect 565759 403348 565771 403382
rect 565805 403348 565817 403382
rect 565759 403307 565817 403348
rect 560555 358948 560613 358989
rect 560555 358914 560567 358948
rect 560601 358914 560613 358948
rect 560555 358880 560613 358914
rect 560555 358846 560567 358880
rect 560601 358846 560613 358880
rect 560555 358812 560613 358846
rect 560555 358778 560567 358812
rect 560601 358778 560613 358812
rect 560555 358744 560613 358778
rect 560555 358710 560567 358744
rect 560601 358710 560613 358744
rect 560555 358676 560613 358710
rect 560555 358642 560567 358676
rect 560601 358642 560613 358676
rect 560555 358608 560613 358642
rect 560555 358574 560567 358608
rect 560601 358574 560613 358608
rect 560555 358540 560613 358574
rect 560555 358506 560567 358540
rect 560601 358506 560613 358540
rect 560555 358472 560613 358506
rect 560555 358438 560567 358472
rect 560601 358438 560613 358472
rect 560555 358404 560613 358438
rect 560555 358370 560567 358404
rect 560601 358370 560613 358404
rect 560555 358336 560613 358370
rect 560555 358302 560567 358336
rect 560601 358302 560613 358336
rect 560555 358268 560613 358302
rect 560555 358234 560567 358268
rect 560601 358234 560613 358268
rect 560555 358200 560613 358234
rect 560555 358166 560567 358200
rect 560601 358166 560613 358200
rect 560555 358132 560613 358166
rect 560555 358098 560567 358132
rect 560601 358098 560613 358132
rect 560555 358064 560613 358098
rect 560555 358030 560567 358064
rect 560601 358030 560613 358064
rect 560555 357989 560613 358030
rect 560813 358948 560871 358989
rect 560813 358914 560825 358948
rect 560859 358914 560871 358948
rect 560813 358880 560871 358914
rect 560813 358846 560825 358880
rect 560859 358846 560871 358880
rect 560813 358812 560871 358846
rect 560813 358778 560825 358812
rect 560859 358778 560871 358812
rect 560813 358744 560871 358778
rect 560813 358710 560825 358744
rect 560859 358710 560871 358744
rect 560813 358676 560871 358710
rect 560813 358642 560825 358676
rect 560859 358642 560871 358676
rect 560813 358608 560871 358642
rect 560813 358574 560825 358608
rect 560859 358574 560871 358608
rect 560813 358540 560871 358574
rect 560813 358506 560825 358540
rect 560859 358506 560871 358540
rect 560813 358472 560871 358506
rect 560813 358438 560825 358472
rect 560859 358438 560871 358472
rect 560813 358404 560871 358438
rect 560813 358370 560825 358404
rect 560859 358370 560871 358404
rect 560813 358336 560871 358370
rect 560813 358302 560825 358336
rect 560859 358302 560871 358336
rect 560813 358268 560871 358302
rect 560813 358234 560825 358268
rect 560859 358234 560871 358268
rect 560813 358200 560871 358234
rect 560813 358166 560825 358200
rect 560859 358166 560871 358200
rect 560813 358132 560871 358166
rect 560813 358098 560825 358132
rect 560859 358098 560871 358132
rect 560813 358064 560871 358098
rect 560813 358030 560825 358064
rect 560859 358030 560871 358064
rect 560813 357989 560871 358030
rect 561071 358948 561129 358989
rect 561071 358914 561083 358948
rect 561117 358914 561129 358948
rect 561071 358880 561129 358914
rect 561071 358846 561083 358880
rect 561117 358846 561129 358880
rect 561071 358812 561129 358846
rect 561071 358778 561083 358812
rect 561117 358778 561129 358812
rect 561071 358744 561129 358778
rect 561071 358710 561083 358744
rect 561117 358710 561129 358744
rect 561071 358676 561129 358710
rect 561071 358642 561083 358676
rect 561117 358642 561129 358676
rect 561071 358608 561129 358642
rect 561071 358574 561083 358608
rect 561117 358574 561129 358608
rect 561071 358540 561129 358574
rect 561071 358506 561083 358540
rect 561117 358506 561129 358540
rect 561071 358472 561129 358506
rect 561071 358438 561083 358472
rect 561117 358438 561129 358472
rect 561071 358404 561129 358438
rect 561071 358370 561083 358404
rect 561117 358370 561129 358404
rect 561071 358336 561129 358370
rect 561071 358302 561083 358336
rect 561117 358302 561129 358336
rect 561071 358268 561129 358302
rect 561071 358234 561083 358268
rect 561117 358234 561129 358268
rect 561071 358200 561129 358234
rect 561071 358166 561083 358200
rect 561117 358166 561129 358200
rect 561071 358132 561129 358166
rect 561071 358098 561083 358132
rect 561117 358098 561129 358132
rect 561071 358064 561129 358098
rect 561071 358030 561083 358064
rect 561117 358030 561129 358064
rect 561071 357989 561129 358030
rect 561329 358948 561387 358989
rect 561329 358914 561341 358948
rect 561375 358914 561387 358948
rect 561329 358880 561387 358914
rect 561329 358846 561341 358880
rect 561375 358846 561387 358880
rect 561329 358812 561387 358846
rect 561329 358778 561341 358812
rect 561375 358778 561387 358812
rect 561329 358744 561387 358778
rect 561329 358710 561341 358744
rect 561375 358710 561387 358744
rect 561329 358676 561387 358710
rect 561329 358642 561341 358676
rect 561375 358642 561387 358676
rect 561329 358608 561387 358642
rect 561329 358574 561341 358608
rect 561375 358574 561387 358608
rect 561329 358540 561387 358574
rect 561329 358506 561341 358540
rect 561375 358506 561387 358540
rect 561329 358472 561387 358506
rect 561329 358438 561341 358472
rect 561375 358438 561387 358472
rect 561329 358404 561387 358438
rect 561329 358370 561341 358404
rect 561375 358370 561387 358404
rect 561329 358336 561387 358370
rect 561329 358302 561341 358336
rect 561375 358302 561387 358336
rect 561329 358268 561387 358302
rect 561329 358234 561341 358268
rect 561375 358234 561387 358268
rect 561329 358200 561387 358234
rect 561329 358166 561341 358200
rect 561375 358166 561387 358200
rect 561329 358132 561387 358166
rect 561329 358098 561341 358132
rect 561375 358098 561387 358132
rect 561329 358064 561387 358098
rect 561329 358030 561341 358064
rect 561375 358030 561387 358064
rect 561329 357989 561387 358030
rect 561587 358948 561645 358989
rect 561587 358914 561599 358948
rect 561633 358914 561645 358948
rect 561587 358880 561645 358914
rect 561587 358846 561599 358880
rect 561633 358846 561645 358880
rect 561587 358812 561645 358846
rect 561587 358778 561599 358812
rect 561633 358778 561645 358812
rect 561587 358744 561645 358778
rect 561587 358710 561599 358744
rect 561633 358710 561645 358744
rect 561587 358676 561645 358710
rect 561587 358642 561599 358676
rect 561633 358642 561645 358676
rect 561587 358608 561645 358642
rect 561587 358574 561599 358608
rect 561633 358574 561645 358608
rect 561587 358540 561645 358574
rect 561587 358506 561599 358540
rect 561633 358506 561645 358540
rect 561587 358472 561645 358506
rect 561587 358438 561599 358472
rect 561633 358438 561645 358472
rect 561587 358404 561645 358438
rect 561587 358370 561599 358404
rect 561633 358370 561645 358404
rect 561587 358336 561645 358370
rect 561587 358302 561599 358336
rect 561633 358302 561645 358336
rect 561587 358268 561645 358302
rect 561587 358234 561599 358268
rect 561633 358234 561645 358268
rect 561587 358200 561645 358234
rect 561587 358166 561599 358200
rect 561633 358166 561645 358200
rect 561587 358132 561645 358166
rect 561587 358098 561599 358132
rect 561633 358098 561645 358132
rect 561587 358064 561645 358098
rect 561587 358030 561599 358064
rect 561633 358030 561645 358064
rect 561587 357989 561645 358030
rect 561845 358948 561903 358989
rect 561845 358914 561857 358948
rect 561891 358914 561903 358948
rect 561845 358880 561903 358914
rect 561845 358846 561857 358880
rect 561891 358846 561903 358880
rect 561845 358812 561903 358846
rect 561845 358778 561857 358812
rect 561891 358778 561903 358812
rect 561845 358744 561903 358778
rect 561845 358710 561857 358744
rect 561891 358710 561903 358744
rect 561845 358676 561903 358710
rect 561845 358642 561857 358676
rect 561891 358642 561903 358676
rect 561845 358608 561903 358642
rect 561845 358574 561857 358608
rect 561891 358574 561903 358608
rect 561845 358540 561903 358574
rect 561845 358506 561857 358540
rect 561891 358506 561903 358540
rect 561845 358472 561903 358506
rect 561845 358438 561857 358472
rect 561891 358438 561903 358472
rect 561845 358404 561903 358438
rect 561845 358370 561857 358404
rect 561891 358370 561903 358404
rect 561845 358336 561903 358370
rect 561845 358302 561857 358336
rect 561891 358302 561903 358336
rect 561845 358268 561903 358302
rect 561845 358234 561857 358268
rect 561891 358234 561903 358268
rect 561845 358200 561903 358234
rect 561845 358166 561857 358200
rect 561891 358166 561903 358200
rect 561845 358132 561903 358166
rect 561845 358098 561857 358132
rect 561891 358098 561903 358132
rect 561845 358064 561903 358098
rect 561845 358030 561857 358064
rect 561891 358030 561903 358064
rect 561845 357989 561903 358030
rect 562103 358948 562161 358989
rect 562103 358914 562115 358948
rect 562149 358914 562161 358948
rect 562103 358880 562161 358914
rect 562103 358846 562115 358880
rect 562149 358846 562161 358880
rect 562103 358812 562161 358846
rect 562103 358778 562115 358812
rect 562149 358778 562161 358812
rect 562103 358744 562161 358778
rect 562103 358710 562115 358744
rect 562149 358710 562161 358744
rect 562103 358676 562161 358710
rect 562103 358642 562115 358676
rect 562149 358642 562161 358676
rect 562103 358608 562161 358642
rect 562103 358574 562115 358608
rect 562149 358574 562161 358608
rect 562103 358540 562161 358574
rect 562103 358506 562115 358540
rect 562149 358506 562161 358540
rect 562103 358472 562161 358506
rect 562103 358438 562115 358472
rect 562149 358438 562161 358472
rect 562103 358404 562161 358438
rect 562103 358370 562115 358404
rect 562149 358370 562161 358404
rect 562103 358336 562161 358370
rect 562103 358302 562115 358336
rect 562149 358302 562161 358336
rect 562103 358268 562161 358302
rect 562103 358234 562115 358268
rect 562149 358234 562161 358268
rect 562103 358200 562161 358234
rect 562103 358166 562115 358200
rect 562149 358166 562161 358200
rect 562103 358132 562161 358166
rect 562103 358098 562115 358132
rect 562149 358098 562161 358132
rect 562103 358064 562161 358098
rect 562103 358030 562115 358064
rect 562149 358030 562161 358064
rect 562103 357989 562161 358030
rect 562361 358948 562419 358989
rect 562361 358914 562373 358948
rect 562407 358914 562419 358948
rect 562361 358880 562419 358914
rect 562361 358846 562373 358880
rect 562407 358846 562419 358880
rect 562361 358812 562419 358846
rect 562361 358778 562373 358812
rect 562407 358778 562419 358812
rect 562361 358744 562419 358778
rect 562361 358710 562373 358744
rect 562407 358710 562419 358744
rect 562361 358676 562419 358710
rect 562361 358642 562373 358676
rect 562407 358642 562419 358676
rect 562361 358608 562419 358642
rect 562361 358574 562373 358608
rect 562407 358574 562419 358608
rect 562361 358540 562419 358574
rect 562361 358506 562373 358540
rect 562407 358506 562419 358540
rect 562361 358472 562419 358506
rect 562361 358438 562373 358472
rect 562407 358438 562419 358472
rect 562361 358404 562419 358438
rect 562361 358370 562373 358404
rect 562407 358370 562419 358404
rect 562361 358336 562419 358370
rect 562361 358302 562373 358336
rect 562407 358302 562419 358336
rect 562361 358268 562419 358302
rect 562361 358234 562373 358268
rect 562407 358234 562419 358268
rect 562361 358200 562419 358234
rect 562361 358166 562373 358200
rect 562407 358166 562419 358200
rect 562361 358132 562419 358166
rect 562361 358098 562373 358132
rect 562407 358098 562419 358132
rect 562361 358064 562419 358098
rect 562361 358030 562373 358064
rect 562407 358030 562419 358064
rect 562361 357989 562419 358030
rect 562619 358948 562677 358989
rect 562619 358914 562631 358948
rect 562665 358914 562677 358948
rect 562619 358880 562677 358914
rect 562619 358846 562631 358880
rect 562665 358846 562677 358880
rect 562619 358812 562677 358846
rect 562619 358778 562631 358812
rect 562665 358778 562677 358812
rect 562619 358744 562677 358778
rect 562619 358710 562631 358744
rect 562665 358710 562677 358744
rect 562619 358676 562677 358710
rect 562619 358642 562631 358676
rect 562665 358642 562677 358676
rect 562619 358608 562677 358642
rect 562619 358574 562631 358608
rect 562665 358574 562677 358608
rect 562619 358540 562677 358574
rect 562619 358506 562631 358540
rect 562665 358506 562677 358540
rect 562619 358472 562677 358506
rect 562619 358438 562631 358472
rect 562665 358438 562677 358472
rect 562619 358404 562677 358438
rect 562619 358370 562631 358404
rect 562665 358370 562677 358404
rect 562619 358336 562677 358370
rect 562619 358302 562631 358336
rect 562665 358302 562677 358336
rect 562619 358268 562677 358302
rect 562619 358234 562631 358268
rect 562665 358234 562677 358268
rect 562619 358200 562677 358234
rect 562619 358166 562631 358200
rect 562665 358166 562677 358200
rect 562619 358132 562677 358166
rect 562619 358098 562631 358132
rect 562665 358098 562677 358132
rect 562619 358064 562677 358098
rect 562619 358030 562631 358064
rect 562665 358030 562677 358064
rect 562619 357989 562677 358030
rect 562877 358948 562935 358989
rect 562877 358914 562889 358948
rect 562923 358914 562935 358948
rect 562877 358880 562935 358914
rect 562877 358846 562889 358880
rect 562923 358846 562935 358880
rect 562877 358812 562935 358846
rect 562877 358778 562889 358812
rect 562923 358778 562935 358812
rect 562877 358744 562935 358778
rect 562877 358710 562889 358744
rect 562923 358710 562935 358744
rect 562877 358676 562935 358710
rect 562877 358642 562889 358676
rect 562923 358642 562935 358676
rect 562877 358608 562935 358642
rect 562877 358574 562889 358608
rect 562923 358574 562935 358608
rect 562877 358540 562935 358574
rect 562877 358506 562889 358540
rect 562923 358506 562935 358540
rect 562877 358472 562935 358506
rect 562877 358438 562889 358472
rect 562923 358438 562935 358472
rect 562877 358404 562935 358438
rect 562877 358370 562889 358404
rect 562923 358370 562935 358404
rect 562877 358336 562935 358370
rect 562877 358302 562889 358336
rect 562923 358302 562935 358336
rect 562877 358268 562935 358302
rect 562877 358234 562889 358268
rect 562923 358234 562935 358268
rect 562877 358200 562935 358234
rect 562877 358166 562889 358200
rect 562923 358166 562935 358200
rect 562877 358132 562935 358166
rect 562877 358098 562889 358132
rect 562923 358098 562935 358132
rect 562877 358064 562935 358098
rect 562877 358030 562889 358064
rect 562923 358030 562935 358064
rect 562877 357989 562935 358030
rect 563135 358948 563193 358989
rect 563135 358914 563147 358948
rect 563181 358914 563193 358948
rect 563135 358880 563193 358914
rect 563135 358846 563147 358880
rect 563181 358846 563193 358880
rect 563135 358812 563193 358846
rect 563135 358778 563147 358812
rect 563181 358778 563193 358812
rect 563135 358744 563193 358778
rect 563135 358710 563147 358744
rect 563181 358710 563193 358744
rect 563135 358676 563193 358710
rect 563135 358642 563147 358676
rect 563181 358642 563193 358676
rect 563135 358608 563193 358642
rect 563135 358574 563147 358608
rect 563181 358574 563193 358608
rect 563135 358540 563193 358574
rect 563135 358506 563147 358540
rect 563181 358506 563193 358540
rect 563135 358472 563193 358506
rect 563135 358438 563147 358472
rect 563181 358438 563193 358472
rect 563135 358404 563193 358438
rect 563135 358370 563147 358404
rect 563181 358370 563193 358404
rect 563135 358336 563193 358370
rect 563135 358302 563147 358336
rect 563181 358302 563193 358336
rect 563135 358268 563193 358302
rect 563135 358234 563147 358268
rect 563181 358234 563193 358268
rect 563135 358200 563193 358234
rect 563135 358166 563147 358200
rect 563181 358166 563193 358200
rect 563135 358132 563193 358166
rect 563135 358098 563147 358132
rect 563181 358098 563193 358132
rect 563135 358064 563193 358098
rect 563135 358030 563147 358064
rect 563181 358030 563193 358064
rect 563135 357989 563193 358030
rect 563393 358948 563451 358989
rect 563393 358914 563405 358948
rect 563439 358914 563451 358948
rect 563393 358880 563451 358914
rect 563393 358846 563405 358880
rect 563439 358846 563451 358880
rect 563393 358812 563451 358846
rect 563393 358778 563405 358812
rect 563439 358778 563451 358812
rect 563393 358744 563451 358778
rect 563393 358710 563405 358744
rect 563439 358710 563451 358744
rect 563393 358676 563451 358710
rect 563393 358642 563405 358676
rect 563439 358642 563451 358676
rect 563393 358608 563451 358642
rect 563393 358574 563405 358608
rect 563439 358574 563451 358608
rect 563393 358540 563451 358574
rect 563393 358506 563405 358540
rect 563439 358506 563451 358540
rect 563393 358472 563451 358506
rect 563393 358438 563405 358472
rect 563439 358438 563451 358472
rect 563393 358404 563451 358438
rect 563393 358370 563405 358404
rect 563439 358370 563451 358404
rect 563393 358336 563451 358370
rect 563393 358302 563405 358336
rect 563439 358302 563451 358336
rect 563393 358268 563451 358302
rect 563393 358234 563405 358268
rect 563439 358234 563451 358268
rect 563393 358200 563451 358234
rect 563393 358166 563405 358200
rect 563439 358166 563451 358200
rect 563393 358132 563451 358166
rect 563393 358098 563405 358132
rect 563439 358098 563451 358132
rect 563393 358064 563451 358098
rect 563393 358030 563405 358064
rect 563439 358030 563451 358064
rect 563393 357989 563451 358030
rect 563651 358948 563709 358989
rect 563651 358914 563663 358948
rect 563697 358914 563709 358948
rect 563651 358880 563709 358914
rect 563651 358846 563663 358880
rect 563697 358846 563709 358880
rect 563651 358812 563709 358846
rect 563651 358778 563663 358812
rect 563697 358778 563709 358812
rect 563651 358744 563709 358778
rect 563651 358710 563663 358744
rect 563697 358710 563709 358744
rect 563651 358676 563709 358710
rect 563651 358642 563663 358676
rect 563697 358642 563709 358676
rect 563651 358608 563709 358642
rect 563651 358574 563663 358608
rect 563697 358574 563709 358608
rect 563651 358540 563709 358574
rect 563651 358506 563663 358540
rect 563697 358506 563709 358540
rect 563651 358472 563709 358506
rect 563651 358438 563663 358472
rect 563697 358438 563709 358472
rect 563651 358404 563709 358438
rect 563651 358370 563663 358404
rect 563697 358370 563709 358404
rect 563651 358336 563709 358370
rect 563651 358302 563663 358336
rect 563697 358302 563709 358336
rect 563651 358268 563709 358302
rect 563651 358234 563663 358268
rect 563697 358234 563709 358268
rect 563651 358200 563709 358234
rect 563651 358166 563663 358200
rect 563697 358166 563709 358200
rect 563651 358132 563709 358166
rect 563651 358098 563663 358132
rect 563697 358098 563709 358132
rect 563651 358064 563709 358098
rect 563651 358030 563663 358064
rect 563697 358030 563709 358064
rect 563651 357989 563709 358030
rect 563909 358948 563967 358989
rect 563909 358914 563921 358948
rect 563955 358914 563967 358948
rect 563909 358880 563967 358914
rect 563909 358846 563921 358880
rect 563955 358846 563967 358880
rect 563909 358812 563967 358846
rect 563909 358778 563921 358812
rect 563955 358778 563967 358812
rect 563909 358744 563967 358778
rect 563909 358710 563921 358744
rect 563955 358710 563967 358744
rect 563909 358676 563967 358710
rect 563909 358642 563921 358676
rect 563955 358642 563967 358676
rect 563909 358608 563967 358642
rect 563909 358574 563921 358608
rect 563955 358574 563967 358608
rect 563909 358540 563967 358574
rect 563909 358506 563921 358540
rect 563955 358506 563967 358540
rect 563909 358472 563967 358506
rect 563909 358438 563921 358472
rect 563955 358438 563967 358472
rect 563909 358404 563967 358438
rect 563909 358370 563921 358404
rect 563955 358370 563967 358404
rect 563909 358336 563967 358370
rect 563909 358302 563921 358336
rect 563955 358302 563967 358336
rect 563909 358268 563967 358302
rect 563909 358234 563921 358268
rect 563955 358234 563967 358268
rect 563909 358200 563967 358234
rect 563909 358166 563921 358200
rect 563955 358166 563967 358200
rect 563909 358132 563967 358166
rect 563909 358098 563921 358132
rect 563955 358098 563967 358132
rect 563909 358064 563967 358098
rect 563909 358030 563921 358064
rect 563955 358030 563967 358064
rect 563909 357989 563967 358030
rect 564167 358948 564225 358989
rect 564167 358914 564179 358948
rect 564213 358914 564225 358948
rect 564167 358880 564225 358914
rect 564167 358846 564179 358880
rect 564213 358846 564225 358880
rect 564167 358812 564225 358846
rect 564167 358778 564179 358812
rect 564213 358778 564225 358812
rect 564167 358744 564225 358778
rect 564167 358710 564179 358744
rect 564213 358710 564225 358744
rect 564167 358676 564225 358710
rect 564167 358642 564179 358676
rect 564213 358642 564225 358676
rect 564167 358608 564225 358642
rect 564167 358574 564179 358608
rect 564213 358574 564225 358608
rect 564167 358540 564225 358574
rect 564167 358506 564179 358540
rect 564213 358506 564225 358540
rect 564167 358472 564225 358506
rect 564167 358438 564179 358472
rect 564213 358438 564225 358472
rect 564167 358404 564225 358438
rect 564167 358370 564179 358404
rect 564213 358370 564225 358404
rect 564167 358336 564225 358370
rect 564167 358302 564179 358336
rect 564213 358302 564225 358336
rect 564167 358268 564225 358302
rect 564167 358234 564179 358268
rect 564213 358234 564225 358268
rect 564167 358200 564225 358234
rect 564167 358166 564179 358200
rect 564213 358166 564225 358200
rect 564167 358132 564225 358166
rect 564167 358098 564179 358132
rect 564213 358098 564225 358132
rect 564167 358064 564225 358098
rect 564167 358030 564179 358064
rect 564213 358030 564225 358064
rect 564167 357989 564225 358030
rect 564425 358948 564483 358989
rect 564425 358914 564437 358948
rect 564471 358914 564483 358948
rect 564425 358880 564483 358914
rect 564425 358846 564437 358880
rect 564471 358846 564483 358880
rect 564425 358812 564483 358846
rect 564425 358778 564437 358812
rect 564471 358778 564483 358812
rect 564425 358744 564483 358778
rect 564425 358710 564437 358744
rect 564471 358710 564483 358744
rect 564425 358676 564483 358710
rect 564425 358642 564437 358676
rect 564471 358642 564483 358676
rect 564425 358608 564483 358642
rect 564425 358574 564437 358608
rect 564471 358574 564483 358608
rect 564425 358540 564483 358574
rect 564425 358506 564437 358540
rect 564471 358506 564483 358540
rect 564425 358472 564483 358506
rect 564425 358438 564437 358472
rect 564471 358438 564483 358472
rect 564425 358404 564483 358438
rect 564425 358370 564437 358404
rect 564471 358370 564483 358404
rect 564425 358336 564483 358370
rect 564425 358302 564437 358336
rect 564471 358302 564483 358336
rect 564425 358268 564483 358302
rect 564425 358234 564437 358268
rect 564471 358234 564483 358268
rect 564425 358200 564483 358234
rect 564425 358166 564437 358200
rect 564471 358166 564483 358200
rect 564425 358132 564483 358166
rect 564425 358098 564437 358132
rect 564471 358098 564483 358132
rect 564425 358064 564483 358098
rect 564425 358030 564437 358064
rect 564471 358030 564483 358064
rect 564425 357989 564483 358030
rect 564683 358948 564741 358989
rect 564683 358914 564695 358948
rect 564729 358914 564741 358948
rect 564683 358880 564741 358914
rect 564683 358846 564695 358880
rect 564729 358846 564741 358880
rect 564683 358812 564741 358846
rect 564683 358778 564695 358812
rect 564729 358778 564741 358812
rect 564683 358744 564741 358778
rect 564683 358710 564695 358744
rect 564729 358710 564741 358744
rect 564683 358676 564741 358710
rect 564683 358642 564695 358676
rect 564729 358642 564741 358676
rect 564683 358608 564741 358642
rect 564683 358574 564695 358608
rect 564729 358574 564741 358608
rect 564683 358540 564741 358574
rect 564683 358506 564695 358540
rect 564729 358506 564741 358540
rect 564683 358472 564741 358506
rect 564683 358438 564695 358472
rect 564729 358438 564741 358472
rect 564683 358404 564741 358438
rect 564683 358370 564695 358404
rect 564729 358370 564741 358404
rect 564683 358336 564741 358370
rect 564683 358302 564695 358336
rect 564729 358302 564741 358336
rect 564683 358268 564741 358302
rect 564683 358234 564695 358268
rect 564729 358234 564741 358268
rect 564683 358200 564741 358234
rect 564683 358166 564695 358200
rect 564729 358166 564741 358200
rect 564683 358132 564741 358166
rect 564683 358098 564695 358132
rect 564729 358098 564741 358132
rect 564683 358064 564741 358098
rect 564683 358030 564695 358064
rect 564729 358030 564741 358064
rect 564683 357989 564741 358030
rect 564941 358948 564999 358989
rect 564941 358914 564953 358948
rect 564987 358914 564999 358948
rect 564941 358880 564999 358914
rect 564941 358846 564953 358880
rect 564987 358846 564999 358880
rect 564941 358812 564999 358846
rect 564941 358778 564953 358812
rect 564987 358778 564999 358812
rect 564941 358744 564999 358778
rect 564941 358710 564953 358744
rect 564987 358710 564999 358744
rect 564941 358676 564999 358710
rect 564941 358642 564953 358676
rect 564987 358642 564999 358676
rect 564941 358608 564999 358642
rect 564941 358574 564953 358608
rect 564987 358574 564999 358608
rect 564941 358540 564999 358574
rect 564941 358506 564953 358540
rect 564987 358506 564999 358540
rect 564941 358472 564999 358506
rect 564941 358438 564953 358472
rect 564987 358438 564999 358472
rect 564941 358404 564999 358438
rect 564941 358370 564953 358404
rect 564987 358370 564999 358404
rect 564941 358336 564999 358370
rect 564941 358302 564953 358336
rect 564987 358302 564999 358336
rect 564941 358268 564999 358302
rect 564941 358234 564953 358268
rect 564987 358234 564999 358268
rect 564941 358200 564999 358234
rect 564941 358166 564953 358200
rect 564987 358166 564999 358200
rect 564941 358132 564999 358166
rect 564941 358098 564953 358132
rect 564987 358098 564999 358132
rect 564941 358064 564999 358098
rect 564941 358030 564953 358064
rect 564987 358030 564999 358064
rect 564941 357989 564999 358030
rect 565199 358948 565257 358989
rect 565199 358914 565211 358948
rect 565245 358914 565257 358948
rect 565199 358880 565257 358914
rect 565199 358846 565211 358880
rect 565245 358846 565257 358880
rect 565199 358812 565257 358846
rect 565199 358778 565211 358812
rect 565245 358778 565257 358812
rect 565199 358744 565257 358778
rect 565199 358710 565211 358744
rect 565245 358710 565257 358744
rect 565199 358676 565257 358710
rect 565199 358642 565211 358676
rect 565245 358642 565257 358676
rect 565199 358608 565257 358642
rect 565199 358574 565211 358608
rect 565245 358574 565257 358608
rect 565199 358540 565257 358574
rect 565199 358506 565211 358540
rect 565245 358506 565257 358540
rect 565199 358472 565257 358506
rect 565199 358438 565211 358472
rect 565245 358438 565257 358472
rect 565199 358404 565257 358438
rect 565199 358370 565211 358404
rect 565245 358370 565257 358404
rect 565199 358336 565257 358370
rect 565199 358302 565211 358336
rect 565245 358302 565257 358336
rect 565199 358268 565257 358302
rect 565199 358234 565211 358268
rect 565245 358234 565257 358268
rect 565199 358200 565257 358234
rect 565199 358166 565211 358200
rect 565245 358166 565257 358200
rect 565199 358132 565257 358166
rect 565199 358098 565211 358132
rect 565245 358098 565257 358132
rect 565199 358064 565257 358098
rect 565199 358030 565211 358064
rect 565245 358030 565257 358064
rect 565199 357989 565257 358030
rect 565457 358948 565515 358989
rect 565457 358914 565469 358948
rect 565503 358914 565515 358948
rect 565457 358880 565515 358914
rect 565457 358846 565469 358880
rect 565503 358846 565515 358880
rect 565457 358812 565515 358846
rect 565457 358778 565469 358812
rect 565503 358778 565515 358812
rect 565457 358744 565515 358778
rect 565457 358710 565469 358744
rect 565503 358710 565515 358744
rect 565457 358676 565515 358710
rect 565457 358642 565469 358676
rect 565503 358642 565515 358676
rect 565457 358608 565515 358642
rect 565457 358574 565469 358608
rect 565503 358574 565515 358608
rect 565457 358540 565515 358574
rect 565457 358506 565469 358540
rect 565503 358506 565515 358540
rect 565457 358472 565515 358506
rect 565457 358438 565469 358472
rect 565503 358438 565515 358472
rect 565457 358404 565515 358438
rect 565457 358370 565469 358404
rect 565503 358370 565515 358404
rect 565457 358336 565515 358370
rect 565457 358302 565469 358336
rect 565503 358302 565515 358336
rect 565457 358268 565515 358302
rect 565457 358234 565469 358268
rect 565503 358234 565515 358268
rect 565457 358200 565515 358234
rect 565457 358166 565469 358200
rect 565503 358166 565515 358200
rect 565457 358132 565515 358166
rect 565457 358098 565469 358132
rect 565503 358098 565515 358132
rect 565457 358064 565515 358098
rect 565457 358030 565469 358064
rect 565503 358030 565515 358064
rect 565457 357989 565515 358030
rect 565715 358948 565773 358989
rect 565715 358914 565727 358948
rect 565761 358914 565773 358948
rect 565715 358880 565773 358914
rect 565715 358846 565727 358880
rect 565761 358846 565773 358880
rect 565715 358812 565773 358846
rect 565715 358778 565727 358812
rect 565761 358778 565773 358812
rect 565715 358744 565773 358778
rect 565715 358710 565727 358744
rect 565761 358710 565773 358744
rect 565715 358676 565773 358710
rect 565715 358642 565727 358676
rect 565761 358642 565773 358676
rect 565715 358608 565773 358642
rect 565715 358574 565727 358608
rect 565761 358574 565773 358608
rect 565715 358540 565773 358574
rect 565715 358506 565727 358540
rect 565761 358506 565773 358540
rect 565715 358472 565773 358506
rect 565715 358438 565727 358472
rect 565761 358438 565773 358472
rect 565715 358404 565773 358438
rect 565715 358370 565727 358404
rect 565761 358370 565773 358404
rect 565715 358336 565773 358370
rect 565715 358302 565727 358336
rect 565761 358302 565773 358336
rect 565715 358268 565773 358302
rect 565715 358234 565727 358268
rect 565761 358234 565773 358268
rect 565715 358200 565773 358234
rect 565715 358166 565727 358200
rect 565761 358166 565773 358200
rect 565715 358132 565773 358166
rect 565715 358098 565727 358132
rect 565761 358098 565773 358132
rect 565715 358064 565773 358098
rect 565715 358030 565727 358064
rect 565761 358030 565773 358064
rect 565715 357989 565773 358030
rect 560417 312640 560475 312681
rect 560417 312606 560429 312640
rect 560463 312606 560475 312640
rect 560417 312572 560475 312606
rect 560417 312538 560429 312572
rect 560463 312538 560475 312572
rect 560417 312504 560475 312538
rect 560417 312470 560429 312504
rect 560463 312470 560475 312504
rect 560417 312436 560475 312470
rect 560417 312402 560429 312436
rect 560463 312402 560475 312436
rect 560417 312368 560475 312402
rect 560417 312334 560429 312368
rect 560463 312334 560475 312368
rect 560417 312300 560475 312334
rect 560417 312266 560429 312300
rect 560463 312266 560475 312300
rect 560417 312232 560475 312266
rect 560417 312198 560429 312232
rect 560463 312198 560475 312232
rect 560417 312164 560475 312198
rect 560417 312130 560429 312164
rect 560463 312130 560475 312164
rect 560417 312096 560475 312130
rect 560417 312062 560429 312096
rect 560463 312062 560475 312096
rect 560417 312028 560475 312062
rect 560417 311994 560429 312028
rect 560463 311994 560475 312028
rect 560417 311960 560475 311994
rect 560417 311926 560429 311960
rect 560463 311926 560475 311960
rect 560417 311892 560475 311926
rect 560417 311858 560429 311892
rect 560463 311858 560475 311892
rect 560417 311824 560475 311858
rect 560417 311790 560429 311824
rect 560463 311790 560475 311824
rect 560417 311756 560475 311790
rect 560417 311722 560429 311756
rect 560463 311722 560475 311756
rect 560417 311681 560475 311722
rect 560675 312640 560733 312681
rect 560675 312606 560687 312640
rect 560721 312606 560733 312640
rect 560675 312572 560733 312606
rect 560675 312538 560687 312572
rect 560721 312538 560733 312572
rect 560675 312504 560733 312538
rect 560675 312470 560687 312504
rect 560721 312470 560733 312504
rect 560675 312436 560733 312470
rect 560675 312402 560687 312436
rect 560721 312402 560733 312436
rect 560675 312368 560733 312402
rect 560675 312334 560687 312368
rect 560721 312334 560733 312368
rect 560675 312300 560733 312334
rect 560675 312266 560687 312300
rect 560721 312266 560733 312300
rect 560675 312232 560733 312266
rect 560675 312198 560687 312232
rect 560721 312198 560733 312232
rect 560675 312164 560733 312198
rect 560675 312130 560687 312164
rect 560721 312130 560733 312164
rect 560675 312096 560733 312130
rect 560675 312062 560687 312096
rect 560721 312062 560733 312096
rect 560675 312028 560733 312062
rect 560675 311994 560687 312028
rect 560721 311994 560733 312028
rect 560675 311960 560733 311994
rect 560675 311926 560687 311960
rect 560721 311926 560733 311960
rect 560675 311892 560733 311926
rect 560675 311858 560687 311892
rect 560721 311858 560733 311892
rect 560675 311824 560733 311858
rect 560675 311790 560687 311824
rect 560721 311790 560733 311824
rect 560675 311756 560733 311790
rect 560675 311722 560687 311756
rect 560721 311722 560733 311756
rect 560675 311681 560733 311722
rect 560933 312640 560991 312681
rect 560933 312606 560945 312640
rect 560979 312606 560991 312640
rect 560933 312572 560991 312606
rect 560933 312538 560945 312572
rect 560979 312538 560991 312572
rect 560933 312504 560991 312538
rect 560933 312470 560945 312504
rect 560979 312470 560991 312504
rect 560933 312436 560991 312470
rect 560933 312402 560945 312436
rect 560979 312402 560991 312436
rect 560933 312368 560991 312402
rect 560933 312334 560945 312368
rect 560979 312334 560991 312368
rect 560933 312300 560991 312334
rect 560933 312266 560945 312300
rect 560979 312266 560991 312300
rect 560933 312232 560991 312266
rect 560933 312198 560945 312232
rect 560979 312198 560991 312232
rect 560933 312164 560991 312198
rect 560933 312130 560945 312164
rect 560979 312130 560991 312164
rect 560933 312096 560991 312130
rect 560933 312062 560945 312096
rect 560979 312062 560991 312096
rect 560933 312028 560991 312062
rect 560933 311994 560945 312028
rect 560979 311994 560991 312028
rect 560933 311960 560991 311994
rect 560933 311926 560945 311960
rect 560979 311926 560991 311960
rect 560933 311892 560991 311926
rect 560933 311858 560945 311892
rect 560979 311858 560991 311892
rect 560933 311824 560991 311858
rect 560933 311790 560945 311824
rect 560979 311790 560991 311824
rect 560933 311756 560991 311790
rect 560933 311722 560945 311756
rect 560979 311722 560991 311756
rect 560933 311681 560991 311722
rect 561191 312640 561249 312681
rect 561191 312606 561203 312640
rect 561237 312606 561249 312640
rect 561191 312572 561249 312606
rect 561191 312538 561203 312572
rect 561237 312538 561249 312572
rect 561191 312504 561249 312538
rect 561191 312470 561203 312504
rect 561237 312470 561249 312504
rect 561191 312436 561249 312470
rect 561191 312402 561203 312436
rect 561237 312402 561249 312436
rect 561191 312368 561249 312402
rect 561191 312334 561203 312368
rect 561237 312334 561249 312368
rect 561191 312300 561249 312334
rect 561191 312266 561203 312300
rect 561237 312266 561249 312300
rect 561191 312232 561249 312266
rect 561191 312198 561203 312232
rect 561237 312198 561249 312232
rect 561191 312164 561249 312198
rect 561191 312130 561203 312164
rect 561237 312130 561249 312164
rect 561191 312096 561249 312130
rect 561191 312062 561203 312096
rect 561237 312062 561249 312096
rect 561191 312028 561249 312062
rect 561191 311994 561203 312028
rect 561237 311994 561249 312028
rect 561191 311960 561249 311994
rect 561191 311926 561203 311960
rect 561237 311926 561249 311960
rect 561191 311892 561249 311926
rect 561191 311858 561203 311892
rect 561237 311858 561249 311892
rect 561191 311824 561249 311858
rect 561191 311790 561203 311824
rect 561237 311790 561249 311824
rect 561191 311756 561249 311790
rect 561191 311722 561203 311756
rect 561237 311722 561249 311756
rect 561191 311681 561249 311722
rect 561449 312640 561507 312681
rect 561449 312606 561461 312640
rect 561495 312606 561507 312640
rect 561449 312572 561507 312606
rect 561449 312538 561461 312572
rect 561495 312538 561507 312572
rect 561449 312504 561507 312538
rect 561449 312470 561461 312504
rect 561495 312470 561507 312504
rect 561449 312436 561507 312470
rect 561449 312402 561461 312436
rect 561495 312402 561507 312436
rect 561449 312368 561507 312402
rect 561449 312334 561461 312368
rect 561495 312334 561507 312368
rect 561449 312300 561507 312334
rect 561449 312266 561461 312300
rect 561495 312266 561507 312300
rect 561449 312232 561507 312266
rect 561449 312198 561461 312232
rect 561495 312198 561507 312232
rect 561449 312164 561507 312198
rect 561449 312130 561461 312164
rect 561495 312130 561507 312164
rect 561449 312096 561507 312130
rect 561449 312062 561461 312096
rect 561495 312062 561507 312096
rect 561449 312028 561507 312062
rect 561449 311994 561461 312028
rect 561495 311994 561507 312028
rect 561449 311960 561507 311994
rect 561449 311926 561461 311960
rect 561495 311926 561507 311960
rect 561449 311892 561507 311926
rect 561449 311858 561461 311892
rect 561495 311858 561507 311892
rect 561449 311824 561507 311858
rect 561449 311790 561461 311824
rect 561495 311790 561507 311824
rect 561449 311756 561507 311790
rect 561449 311722 561461 311756
rect 561495 311722 561507 311756
rect 561449 311681 561507 311722
rect 561707 312640 561765 312681
rect 561707 312606 561719 312640
rect 561753 312606 561765 312640
rect 561707 312572 561765 312606
rect 561707 312538 561719 312572
rect 561753 312538 561765 312572
rect 561707 312504 561765 312538
rect 561707 312470 561719 312504
rect 561753 312470 561765 312504
rect 561707 312436 561765 312470
rect 561707 312402 561719 312436
rect 561753 312402 561765 312436
rect 561707 312368 561765 312402
rect 561707 312334 561719 312368
rect 561753 312334 561765 312368
rect 561707 312300 561765 312334
rect 561707 312266 561719 312300
rect 561753 312266 561765 312300
rect 561707 312232 561765 312266
rect 561707 312198 561719 312232
rect 561753 312198 561765 312232
rect 561707 312164 561765 312198
rect 561707 312130 561719 312164
rect 561753 312130 561765 312164
rect 561707 312096 561765 312130
rect 561707 312062 561719 312096
rect 561753 312062 561765 312096
rect 561707 312028 561765 312062
rect 561707 311994 561719 312028
rect 561753 311994 561765 312028
rect 561707 311960 561765 311994
rect 561707 311926 561719 311960
rect 561753 311926 561765 311960
rect 561707 311892 561765 311926
rect 561707 311858 561719 311892
rect 561753 311858 561765 311892
rect 561707 311824 561765 311858
rect 561707 311790 561719 311824
rect 561753 311790 561765 311824
rect 561707 311756 561765 311790
rect 561707 311722 561719 311756
rect 561753 311722 561765 311756
rect 561707 311681 561765 311722
rect 561965 312640 562023 312681
rect 561965 312606 561977 312640
rect 562011 312606 562023 312640
rect 561965 312572 562023 312606
rect 561965 312538 561977 312572
rect 562011 312538 562023 312572
rect 561965 312504 562023 312538
rect 561965 312470 561977 312504
rect 562011 312470 562023 312504
rect 561965 312436 562023 312470
rect 561965 312402 561977 312436
rect 562011 312402 562023 312436
rect 561965 312368 562023 312402
rect 561965 312334 561977 312368
rect 562011 312334 562023 312368
rect 561965 312300 562023 312334
rect 561965 312266 561977 312300
rect 562011 312266 562023 312300
rect 561965 312232 562023 312266
rect 561965 312198 561977 312232
rect 562011 312198 562023 312232
rect 561965 312164 562023 312198
rect 561965 312130 561977 312164
rect 562011 312130 562023 312164
rect 561965 312096 562023 312130
rect 561965 312062 561977 312096
rect 562011 312062 562023 312096
rect 561965 312028 562023 312062
rect 561965 311994 561977 312028
rect 562011 311994 562023 312028
rect 561965 311960 562023 311994
rect 561965 311926 561977 311960
rect 562011 311926 562023 311960
rect 561965 311892 562023 311926
rect 561965 311858 561977 311892
rect 562011 311858 562023 311892
rect 561965 311824 562023 311858
rect 561965 311790 561977 311824
rect 562011 311790 562023 311824
rect 561965 311756 562023 311790
rect 561965 311722 561977 311756
rect 562011 311722 562023 311756
rect 561965 311681 562023 311722
rect 562223 312640 562281 312681
rect 562223 312606 562235 312640
rect 562269 312606 562281 312640
rect 562223 312572 562281 312606
rect 562223 312538 562235 312572
rect 562269 312538 562281 312572
rect 562223 312504 562281 312538
rect 562223 312470 562235 312504
rect 562269 312470 562281 312504
rect 562223 312436 562281 312470
rect 562223 312402 562235 312436
rect 562269 312402 562281 312436
rect 562223 312368 562281 312402
rect 562223 312334 562235 312368
rect 562269 312334 562281 312368
rect 562223 312300 562281 312334
rect 562223 312266 562235 312300
rect 562269 312266 562281 312300
rect 562223 312232 562281 312266
rect 562223 312198 562235 312232
rect 562269 312198 562281 312232
rect 562223 312164 562281 312198
rect 562223 312130 562235 312164
rect 562269 312130 562281 312164
rect 562223 312096 562281 312130
rect 562223 312062 562235 312096
rect 562269 312062 562281 312096
rect 562223 312028 562281 312062
rect 562223 311994 562235 312028
rect 562269 311994 562281 312028
rect 562223 311960 562281 311994
rect 562223 311926 562235 311960
rect 562269 311926 562281 311960
rect 562223 311892 562281 311926
rect 562223 311858 562235 311892
rect 562269 311858 562281 311892
rect 562223 311824 562281 311858
rect 562223 311790 562235 311824
rect 562269 311790 562281 311824
rect 562223 311756 562281 311790
rect 562223 311722 562235 311756
rect 562269 311722 562281 311756
rect 562223 311681 562281 311722
rect 562481 312640 562539 312681
rect 562481 312606 562493 312640
rect 562527 312606 562539 312640
rect 562481 312572 562539 312606
rect 562481 312538 562493 312572
rect 562527 312538 562539 312572
rect 562481 312504 562539 312538
rect 562481 312470 562493 312504
rect 562527 312470 562539 312504
rect 562481 312436 562539 312470
rect 562481 312402 562493 312436
rect 562527 312402 562539 312436
rect 562481 312368 562539 312402
rect 562481 312334 562493 312368
rect 562527 312334 562539 312368
rect 562481 312300 562539 312334
rect 562481 312266 562493 312300
rect 562527 312266 562539 312300
rect 562481 312232 562539 312266
rect 562481 312198 562493 312232
rect 562527 312198 562539 312232
rect 562481 312164 562539 312198
rect 562481 312130 562493 312164
rect 562527 312130 562539 312164
rect 562481 312096 562539 312130
rect 562481 312062 562493 312096
rect 562527 312062 562539 312096
rect 562481 312028 562539 312062
rect 562481 311994 562493 312028
rect 562527 311994 562539 312028
rect 562481 311960 562539 311994
rect 562481 311926 562493 311960
rect 562527 311926 562539 311960
rect 562481 311892 562539 311926
rect 562481 311858 562493 311892
rect 562527 311858 562539 311892
rect 562481 311824 562539 311858
rect 562481 311790 562493 311824
rect 562527 311790 562539 311824
rect 562481 311756 562539 311790
rect 562481 311722 562493 311756
rect 562527 311722 562539 311756
rect 562481 311681 562539 311722
rect 562739 312640 562797 312681
rect 562739 312606 562751 312640
rect 562785 312606 562797 312640
rect 562739 312572 562797 312606
rect 562739 312538 562751 312572
rect 562785 312538 562797 312572
rect 562739 312504 562797 312538
rect 562739 312470 562751 312504
rect 562785 312470 562797 312504
rect 562739 312436 562797 312470
rect 562739 312402 562751 312436
rect 562785 312402 562797 312436
rect 562739 312368 562797 312402
rect 562739 312334 562751 312368
rect 562785 312334 562797 312368
rect 562739 312300 562797 312334
rect 562739 312266 562751 312300
rect 562785 312266 562797 312300
rect 562739 312232 562797 312266
rect 562739 312198 562751 312232
rect 562785 312198 562797 312232
rect 562739 312164 562797 312198
rect 562739 312130 562751 312164
rect 562785 312130 562797 312164
rect 562739 312096 562797 312130
rect 562739 312062 562751 312096
rect 562785 312062 562797 312096
rect 562739 312028 562797 312062
rect 562739 311994 562751 312028
rect 562785 311994 562797 312028
rect 562739 311960 562797 311994
rect 562739 311926 562751 311960
rect 562785 311926 562797 311960
rect 562739 311892 562797 311926
rect 562739 311858 562751 311892
rect 562785 311858 562797 311892
rect 562739 311824 562797 311858
rect 562739 311790 562751 311824
rect 562785 311790 562797 311824
rect 562739 311756 562797 311790
rect 562739 311722 562751 311756
rect 562785 311722 562797 311756
rect 562739 311681 562797 311722
rect 562997 312640 563055 312681
rect 562997 312606 563009 312640
rect 563043 312606 563055 312640
rect 562997 312572 563055 312606
rect 562997 312538 563009 312572
rect 563043 312538 563055 312572
rect 562997 312504 563055 312538
rect 562997 312470 563009 312504
rect 563043 312470 563055 312504
rect 562997 312436 563055 312470
rect 562997 312402 563009 312436
rect 563043 312402 563055 312436
rect 562997 312368 563055 312402
rect 562997 312334 563009 312368
rect 563043 312334 563055 312368
rect 562997 312300 563055 312334
rect 562997 312266 563009 312300
rect 563043 312266 563055 312300
rect 562997 312232 563055 312266
rect 562997 312198 563009 312232
rect 563043 312198 563055 312232
rect 562997 312164 563055 312198
rect 562997 312130 563009 312164
rect 563043 312130 563055 312164
rect 562997 312096 563055 312130
rect 562997 312062 563009 312096
rect 563043 312062 563055 312096
rect 562997 312028 563055 312062
rect 562997 311994 563009 312028
rect 563043 311994 563055 312028
rect 562997 311960 563055 311994
rect 562997 311926 563009 311960
rect 563043 311926 563055 311960
rect 562997 311892 563055 311926
rect 562997 311858 563009 311892
rect 563043 311858 563055 311892
rect 562997 311824 563055 311858
rect 562997 311790 563009 311824
rect 563043 311790 563055 311824
rect 562997 311756 563055 311790
rect 562997 311722 563009 311756
rect 563043 311722 563055 311756
rect 562997 311681 563055 311722
rect 563255 312640 563313 312681
rect 563255 312606 563267 312640
rect 563301 312606 563313 312640
rect 563255 312572 563313 312606
rect 563255 312538 563267 312572
rect 563301 312538 563313 312572
rect 563255 312504 563313 312538
rect 563255 312470 563267 312504
rect 563301 312470 563313 312504
rect 563255 312436 563313 312470
rect 563255 312402 563267 312436
rect 563301 312402 563313 312436
rect 563255 312368 563313 312402
rect 563255 312334 563267 312368
rect 563301 312334 563313 312368
rect 563255 312300 563313 312334
rect 563255 312266 563267 312300
rect 563301 312266 563313 312300
rect 563255 312232 563313 312266
rect 563255 312198 563267 312232
rect 563301 312198 563313 312232
rect 563255 312164 563313 312198
rect 563255 312130 563267 312164
rect 563301 312130 563313 312164
rect 563255 312096 563313 312130
rect 563255 312062 563267 312096
rect 563301 312062 563313 312096
rect 563255 312028 563313 312062
rect 563255 311994 563267 312028
rect 563301 311994 563313 312028
rect 563255 311960 563313 311994
rect 563255 311926 563267 311960
rect 563301 311926 563313 311960
rect 563255 311892 563313 311926
rect 563255 311858 563267 311892
rect 563301 311858 563313 311892
rect 563255 311824 563313 311858
rect 563255 311790 563267 311824
rect 563301 311790 563313 311824
rect 563255 311756 563313 311790
rect 563255 311722 563267 311756
rect 563301 311722 563313 311756
rect 563255 311681 563313 311722
rect 563513 312640 563571 312681
rect 563513 312606 563525 312640
rect 563559 312606 563571 312640
rect 563513 312572 563571 312606
rect 563513 312538 563525 312572
rect 563559 312538 563571 312572
rect 563513 312504 563571 312538
rect 563513 312470 563525 312504
rect 563559 312470 563571 312504
rect 563513 312436 563571 312470
rect 563513 312402 563525 312436
rect 563559 312402 563571 312436
rect 563513 312368 563571 312402
rect 563513 312334 563525 312368
rect 563559 312334 563571 312368
rect 563513 312300 563571 312334
rect 563513 312266 563525 312300
rect 563559 312266 563571 312300
rect 563513 312232 563571 312266
rect 563513 312198 563525 312232
rect 563559 312198 563571 312232
rect 563513 312164 563571 312198
rect 563513 312130 563525 312164
rect 563559 312130 563571 312164
rect 563513 312096 563571 312130
rect 563513 312062 563525 312096
rect 563559 312062 563571 312096
rect 563513 312028 563571 312062
rect 563513 311994 563525 312028
rect 563559 311994 563571 312028
rect 563513 311960 563571 311994
rect 563513 311926 563525 311960
rect 563559 311926 563571 311960
rect 563513 311892 563571 311926
rect 563513 311858 563525 311892
rect 563559 311858 563571 311892
rect 563513 311824 563571 311858
rect 563513 311790 563525 311824
rect 563559 311790 563571 311824
rect 563513 311756 563571 311790
rect 563513 311722 563525 311756
rect 563559 311722 563571 311756
rect 563513 311681 563571 311722
rect 563771 312640 563829 312681
rect 563771 312606 563783 312640
rect 563817 312606 563829 312640
rect 563771 312572 563829 312606
rect 563771 312538 563783 312572
rect 563817 312538 563829 312572
rect 563771 312504 563829 312538
rect 563771 312470 563783 312504
rect 563817 312470 563829 312504
rect 563771 312436 563829 312470
rect 563771 312402 563783 312436
rect 563817 312402 563829 312436
rect 563771 312368 563829 312402
rect 563771 312334 563783 312368
rect 563817 312334 563829 312368
rect 563771 312300 563829 312334
rect 563771 312266 563783 312300
rect 563817 312266 563829 312300
rect 563771 312232 563829 312266
rect 563771 312198 563783 312232
rect 563817 312198 563829 312232
rect 563771 312164 563829 312198
rect 563771 312130 563783 312164
rect 563817 312130 563829 312164
rect 563771 312096 563829 312130
rect 563771 312062 563783 312096
rect 563817 312062 563829 312096
rect 563771 312028 563829 312062
rect 563771 311994 563783 312028
rect 563817 311994 563829 312028
rect 563771 311960 563829 311994
rect 563771 311926 563783 311960
rect 563817 311926 563829 311960
rect 563771 311892 563829 311926
rect 563771 311858 563783 311892
rect 563817 311858 563829 311892
rect 563771 311824 563829 311858
rect 563771 311790 563783 311824
rect 563817 311790 563829 311824
rect 563771 311756 563829 311790
rect 563771 311722 563783 311756
rect 563817 311722 563829 311756
rect 563771 311681 563829 311722
rect 564029 312640 564087 312681
rect 564029 312606 564041 312640
rect 564075 312606 564087 312640
rect 564029 312572 564087 312606
rect 564029 312538 564041 312572
rect 564075 312538 564087 312572
rect 564029 312504 564087 312538
rect 564029 312470 564041 312504
rect 564075 312470 564087 312504
rect 564029 312436 564087 312470
rect 564029 312402 564041 312436
rect 564075 312402 564087 312436
rect 564029 312368 564087 312402
rect 564029 312334 564041 312368
rect 564075 312334 564087 312368
rect 564029 312300 564087 312334
rect 564029 312266 564041 312300
rect 564075 312266 564087 312300
rect 564029 312232 564087 312266
rect 564029 312198 564041 312232
rect 564075 312198 564087 312232
rect 564029 312164 564087 312198
rect 564029 312130 564041 312164
rect 564075 312130 564087 312164
rect 564029 312096 564087 312130
rect 564029 312062 564041 312096
rect 564075 312062 564087 312096
rect 564029 312028 564087 312062
rect 564029 311994 564041 312028
rect 564075 311994 564087 312028
rect 564029 311960 564087 311994
rect 564029 311926 564041 311960
rect 564075 311926 564087 311960
rect 564029 311892 564087 311926
rect 564029 311858 564041 311892
rect 564075 311858 564087 311892
rect 564029 311824 564087 311858
rect 564029 311790 564041 311824
rect 564075 311790 564087 311824
rect 564029 311756 564087 311790
rect 564029 311722 564041 311756
rect 564075 311722 564087 311756
rect 564029 311681 564087 311722
rect 564287 312640 564345 312681
rect 564287 312606 564299 312640
rect 564333 312606 564345 312640
rect 564287 312572 564345 312606
rect 564287 312538 564299 312572
rect 564333 312538 564345 312572
rect 564287 312504 564345 312538
rect 564287 312470 564299 312504
rect 564333 312470 564345 312504
rect 564287 312436 564345 312470
rect 564287 312402 564299 312436
rect 564333 312402 564345 312436
rect 564287 312368 564345 312402
rect 564287 312334 564299 312368
rect 564333 312334 564345 312368
rect 564287 312300 564345 312334
rect 564287 312266 564299 312300
rect 564333 312266 564345 312300
rect 564287 312232 564345 312266
rect 564287 312198 564299 312232
rect 564333 312198 564345 312232
rect 564287 312164 564345 312198
rect 564287 312130 564299 312164
rect 564333 312130 564345 312164
rect 564287 312096 564345 312130
rect 564287 312062 564299 312096
rect 564333 312062 564345 312096
rect 564287 312028 564345 312062
rect 564287 311994 564299 312028
rect 564333 311994 564345 312028
rect 564287 311960 564345 311994
rect 564287 311926 564299 311960
rect 564333 311926 564345 311960
rect 564287 311892 564345 311926
rect 564287 311858 564299 311892
rect 564333 311858 564345 311892
rect 564287 311824 564345 311858
rect 564287 311790 564299 311824
rect 564333 311790 564345 311824
rect 564287 311756 564345 311790
rect 564287 311722 564299 311756
rect 564333 311722 564345 311756
rect 564287 311681 564345 311722
rect 564545 312640 564603 312681
rect 564545 312606 564557 312640
rect 564591 312606 564603 312640
rect 564545 312572 564603 312606
rect 564545 312538 564557 312572
rect 564591 312538 564603 312572
rect 564545 312504 564603 312538
rect 564545 312470 564557 312504
rect 564591 312470 564603 312504
rect 564545 312436 564603 312470
rect 564545 312402 564557 312436
rect 564591 312402 564603 312436
rect 564545 312368 564603 312402
rect 564545 312334 564557 312368
rect 564591 312334 564603 312368
rect 564545 312300 564603 312334
rect 564545 312266 564557 312300
rect 564591 312266 564603 312300
rect 564545 312232 564603 312266
rect 564545 312198 564557 312232
rect 564591 312198 564603 312232
rect 564545 312164 564603 312198
rect 564545 312130 564557 312164
rect 564591 312130 564603 312164
rect 564545 312096 564603 312130
rect 564545 312062 564557 312096
rect 564591 312062 564603 312096
rect 564545 312028 564603 312062
rect 564545 311994 564557 312028
rect 564591 311994 564603 312028
rect 564545 311960 564603 311994
rect 564545 311926 564557 311960
rect 564591 311926 564603 311960
rect 564545 311892 564603 311926
rect 564545 311858 564557 311892
rect 564591 311858 564603 311892
rect 564545 311824 564603 311858
rect 564545 311790 564557 311824
rect 564591 311790 564603 311824
rect 564545 311756 564603 311790
rect 564545 311722 564557 311756
rect 564591 311722 564603 311756
rect 564545 311681 564603 311722
rect 564803 312640 564861 312681
rect 564803 312606 564815 312640
rect 564849 312606 564861 312640
rect 564803 312572 564861 312606
rect 564803 312538 564815 312572
rect 564849 312538 564861 312572
rect 564803 312504 564861 312538
rect 564803 312470 564815 312504
rect 564849 312470 564861 312504
rect 564803 312436 564861 312470
rect 564803 312402 564815 312436
rect 564849 312402 564861 312436
rect 564803 312368 564861 312402
rect 564803 312334 564815 312368
rect 564849 312334 564861 312368
rect 564803 312300 564861 312334
rect 564803 312266 564815 312300
rect 564849 312266 564861 312300
rect 564803 312232 564861 312266
rect 564803 312198 564815 312232
rect 564849 312198 564861 312232
rect 564803 312164 564861 312198
rect 564803 312130 564815 312164
rect 564849 312130 564861 312164
rect 564803 312096 564861 312130
rect 564803 312062 564815 312096
rect 564849 312062 564861 312096
rect 564803 312028 564861 312062
rect 564803 311994 564815 312028
rect 564849 311994 564861 312028
rect 564803 311960 564861 311994
rect 564803 311926 564815 311960
rect 564849 311926 564861 311960
rect 564803 311892 564861 311926
rect 564803 311858 564815 311892
rect 564849 311858 564861 311892
rect 564803 311824 564861 311858
rect 564803 311790 564815 311824
rect 564849 311790 564861 311824
rect 564803 311756 564861 311790
rect 564803 311722 564815 311756
rect 564849 311722 564861 311756
rect 564803 311681 564861 311722
rect 565061 312640 565119 312681
rect 565061 312606 565073 312640
rect 565107 312606 565119 312640
rect 565061 312572 565119 312606
rect 565061 312538 565073 312572
rect 565107 312538 565119 312572
rect 565061 312504 565119 312538
rect 565061 312470 565073 312504
rect 565107 312470 565119 312504
rect 565061 312436 565119 312470
rect 565061 312402 565073 312436
rect 565107 312402 565119 312436
rect 565061 312368 565119 312402
rect 565061 312334 565073 312368
rect 565107 312334 565119 312368
rect 565061 312300 565119 312334
rect 565061 312266 565073 312300
rect 565107 312266 565119 312300
rect 565061 312232 565119 312266
rect 565061 312198 565073 312232
rect 565107 312198 565119 312232
rect 565061 312164 565119 312198
rect 565061 312130 565073 312164
rect 565107 312130 565119 312164
rect 565061 312096 565119 312130
rect 565061 312062 565073 312096
rect 565107 312062 565119 312096
rect 565061 312028 565119 312062
rect 565061 311994 565073 312028
rect 565107 311994 565119 312028
rect 565061 311960 565119 311994
rect 565061 311926 565073 311960
rect 565107 311926 565119 311960
rect 565061 311892 565119 311926
rect 565061 311858 565073 311892
rect 565107 311858 565119 311892
rect 565061 311824 565119 311858
rect 565061 311790 565073 311824
rect 565107 311790 565119 311824
rect 565061 311756 565119 311790
rect 565061 311722 565073 311756
rect 565107 311722 565119 311756
rect 565061 311681 565119 311722
rect 565319 312640 565377 312681
rect 565319 312606 565331 312640
rect 565365 312606 565377 312640
rect 565319 312572 565377 312606
rect 565319 312538 565331 312572
rect 565365 312538 565377 312572
rect 565319 312504 565377 312538
rect 565319 312470 565331 312504
rect 565365 312470 565377 312504
rect 565319 312436 565377 312470
rect 565319 312402 565331 312436
rect 565365 312402 565377 312436
rect 565319 312368 565377 312402
rect 565319 312334 565331 312368
rect 565365 312334 565377 312368
rect 565319 312300 565377 312334
rect 565319 312266 565331 312300
rect 565365 312266 565377 312300
rect 565319 312232 565377 312266
rect 565319 312198 565331 312232
rect 565365 312198 565377 312232
rect 565319 312164 565377 312198
rect 565319 312130 565331 312164
rect 565365 312130 565377 312164
rect 565319 312096 565377 312130
rect 565319 312062 565331 312096
rect 565365 312062 565377 312096
rect 565319 312028 565377 312062
rect 565319 311994 565331 312028
rect 565365 311994 565377 312028
rect 565319 311960 565377 311994
rect 565319 311926 565331 311960
rect 565365 311926 565377 311960
rect 565319 311892 565377 311926
rect 565319 311858 565331 311892
rect 565365 311858 565377 311892
rect 565319 311824 565377 311858
rect 565319 311790 565331 311824
rect 565365 311790 565377 311824
rect 565319 311756 565377 311790
rect 565319 311722 565331 311756
rect 565365 311722 565377 311756
rect 565319 311681 565377 311722
rect 565577 312640 565635 312681
rect 565577 312606 565589 312640
rect 565623 312606 565635 312640
rect 565577 312572 565635 312606
rect 565577 312538 565589 312572
rect 565623 312538 565635 312572
rect 565577 312504 565635 312538
rect 565577 312470 565589 312504
rect 565623 312470 565635 312504
rect 565577 312436 565635 312470
rect 565577 312402 565589 312436
rect 565623 312402 565635 312436
rect 565577 312368 565635 312402
rect 565577 312334 565589 312368
rect 565623 312334 565635 312368
rect 565577 312300 565635 312334
rect 565577 312266 565589 312300
rect 565623 312266 565635 312300
rect 565577 312232 565635 312266
rect 565577 312198 565589 312232
rect 565623 312198 565635 312232
rect 565577 312164 565635 312198
rect 565577 312130 565589 312164
rect 565623 312130 565635 312164
rect 565577 312096 565635 312130
rect 565577 312062 565589 312096
rect 565623 312062 565635 312096
rect 565577 312028 565635 312062
rect 565577 311994 565589 312028
rect 565623 311994 565635 312028
rect 565577 311960 565635 311994
rect 565577 311926 565589 311960
rect 565623 311926 565635 311960
rect 565577 311892 565635 311926
rect 565577 311858 565589 311892
rect 565623 311858 565635 311892
rect 565577 311824 565635 311858
rect 565577 311790 565589 311824
rect 565623 311790 565635 311824
rect 565577 311756 565635 311790
rect 565577 311722 565589 311756
rect 565623 311722 565635 311756
rect 565577 311681 565635 311722
<< pdiff >>
rect 575219 493182 575277 493223
rect 575219 493148 575231 493182
rect 575265 493148 575277 493182
rect 575219 493114 575277 493148
rect 575219 493080 575231 493114
rect 575265 493080 575277 493114
rect 575219 493046 575277 493080
rect 575219 493012 575231 493046
rect 575265 493012 575277 493046
rect 575219 492978 575277 493012
rect 575219 492944 575231 492978
rect 575265 492944 575277 492978
rect 575219 492910 575277 492944
rect 575219 492876 575231 492910
rect 575265 492876 575277 492910
rect 575219 492842 575277 492876
rect 575219 492808 575231 492842
rect 575265 492808 575277 492842
rect 575219 492774 575277 492808
rect 575219 492740 575231 492774
rect 575265 492740 575277 492774
rect 575219 492706 575277 492740
rect 575219 492672 575231 492706
rect 575265 492672 575277 492706
rect 575219 492638 575277 492672
rect 575219 492604 575231 492638
rect 575265 492604 575277 492638
rect 575219 492570 575277 492604
rect 575219 492536 575231 492570
rect 575265 492536 575277 492570
rect 575219 492502 575277 492536
rect 575219 492468 575231 492502
rect 575265 492468 575277 492502
rect 575219 492434 575277 492468
rect 575219 492400 575231 492434
rect 575265 492400 575277 492434
rect 575219 492366 575277 492400
rect 575219 492332 575231 492366
rect 575265 492332 575277 492366
rect 575219 492298 575277 492332
rect 575219 492264 575231 492298
rect 575265 492264 575277 492298
rect 575219 492223 575277 492264
rect 575477 493182 575535 493223
rect 575477 493148 575489 493182
rect 575523 493148 575535 493182
rect 575477 493114 575535 493148
rect 575477 493080 575489 493114
rect 575523 493080 575535 493114
rect 575477 493046 575535 493080
rect 575477 493012 575489 493046
rect 575523 493012 575535 493046
rect 575477 492978 575535 493012
rect 575477 492944 575489 492978
rect 575523 492944 575535 492978
rect 575477 492910 575535 492944
rect 575477 492876 575489 492910
rect 575523 492876 575535 492910
rect 575477 492842 575535 492876
rect 575477 492808 575489 492842
rect 575523 492808 575535 492842
rect 575477 492774 575535 492808
rect 575477 492740 575489 492774
rect 575523 492740 575535 492774
rect 575477 492706 575535 492740
rect 575477 492672 575489 492706
rect 575523 492672 575535 492706
rect 575477 492638 575535 492672
rect 575477 492604 575489 492638
rect 575523 492604 575535 492638
rect 575477 492570 575535 492604
rect 575477 492536 575489 492570
rect 575523 492536 575535 492570
rect 575477 492502 575535 492536
rect 575477 492468 575489 492502
rect 575523 492468 575535 492502
rect 575477 492434 575535 492468
rect 575477 492400 575489 492434
rect 575523 492400 575535 492434
rect 575477 492366 575535 492400
rect 575477 492332 575489 492366
rect 575523 492332 575535 492366
rect 575477 492298 575535 492332
rect 575477 492264 575489 492298
rect 575523 492264 575535 492298
rect 575477 492223 575535 492264
rect 575735 493182 575793 493223
rect 575735 493148 575747 493182
rect 575781 493148 575793 493182
rect 575735 493114 575793 493148
rect 575735 493080 575747 493114
rect 575781 493080 575793 493114
rect 575735 493046 575793 493080
rect 575735 493012 575747 493046
rect 575781 493012 575793 493046
rect 575735 492978 575793 493012
rect 575735 492944 575747 492978
rect 575781 492944 575793 492978
rect 575735 492910 575793 492944
rect 575735 492876 575747 492910
rect 575781 492876 575793 492910
rect 575735 492842 575793 492876
rect 575735 492808 575747 492842
rect 575781 492808 575793 492842
rect 575735 492774 575793 492808
rect 575735 492740 575747 492774
rect 575781 492740 575793 492774
rect 575735 492706 575793 492740
rect 575735 492672 575747 492706
rect 575781 492672 575793 492706
rect 575735 492638 575793 492672
rect 575735 492604 575747 492638
rect 575781 492604 575793 492638
rect 575735 492570 575793 492604
rect 575735 492536 575747 492570
rect 575781 492536 575793 492570
rect 575735 492502 575793 492536
rect 575735 492468 575747 492502
rect 575781 492468 575793 492502
rect 575735 492434 575793 492468
rect 575735 492400 575747 492434
rect 575781 492400 575793 492434
rect 575735 492366 575793 492400
rect 575735 492332 575747 492366
rect 575781 492332 575793 492366
rect 575735 492298 575793 492332
rect 575735 492264 575747 492298
rect 575781 492264 575793 492298
rect 575735 492223 575793 492264
rect 575993 493182 576051 493223
rect 575993 493148 576005 493182
rect 576039 493148 576051 493182
rect 575993 493114 576051 493148
rect 575993 493080 576005 493114
rect 576039 493080 576051 493114
rect 575993 493046 576051 493080
rect 575993 493012 576005 493046
rect 576039 493012 576051 493046
rect 575993 492978 576051 493012
rect 575993 492944 576005 492978
rect 576039 492944 576051 492978
rect 575993 492910 576051 492944
rect 575993 492876 576005 492910
rect 576039 492876 576051 492910
rect 575993 492842 576051 492876
rect 575993 492808 576005 492842
rect 576039 492808 576051 492842
rect 575993 492774 576051 492808
rect 575993 492740 576005 492774
rect 576039 492740 576051 492774
rect 575993 492706 576051 492740
rect 575993 492672 576005 492706
rect 576039 492672 576051 492706
rect 575993 492638 576051 492672
rect 575993 492604 576005 492638
rect 576039 492604 576051 492638
rect 575993 492570 576051 492604
rect 575993 492536 576005 492570
rect 576039 492536 576051 492570
rect 575993 492502 576051 492536
rect 575993 492468 576005 492502
rect 576039 492468 576051 492502
rect 575993 492434 576051 492468
rect 575993 492400 576005 492434
rect 576039 492400 576051 492434
rect 575993 492366 576051 492400
rect 575993 492332 576005 492366
rect 576039 492332 576051 492366
rect 575993 492298 576051 492332
rect 575993 492264 576005 492298
rect 576039 492264 576051 492298
rect 575993 492223 576051 492264
rect 576251 493182 576309 493223
rect 576251 493148 576263 493182
rect 576297 493148 576309 493182
rect 576251 493114 576309 493148
rect 576251 493080 576263 493114
rect 576297 493080 576309 493114
rect 576251 493046 576309 493080
rect 576251 493012 576263 493046
rect 576297 493012 576309 493046
rect 576251 492978 576309 493012
rect 576251 492944 576263 492978
rect 576297 492944 576309 492978
rect 576251 492910 576309 492944
rect 576251 492876 576263 492910
rect 576297 492876 576309 492910
rect 576251 492842 576309 492876
rect 576251 492808 576263 492842
rect 576297 492808 576309 492842
rect 576251 492774 576309 492808
rect 576251 492740 576263 492774
rect 576297 492740 576309 492774
rect 576251 492706 576309 492740
rect 576251 492672 576263 492706
rect 576297 492672 576309 492706
rect 576251 492638 576309 492672
rect 576251 492604 576263 492638
rect 576297 492604 576309 492638
rect 576251 492570 576309 492604
rect 576251 492536 576263 492570
rect 576297 492536 576309 492570
rect 576251 492502 576309 492536
rect 576251 492468 576263 492502
rect 576297 492468 576309 492502
rect 576251 492434 576309 492468
rect 576251 492400 576263 492434
rect 576297 492400 576309 492434
rect 576251 492366 576309 492400
rect 576251 492332 576263 492366
rect 576297 492332 576309 492366
rect 576251 492298 576309 492332
rect 576251 492264 576263 492298
rect 576297 492264 576309 492298
rect 576251 492223 576309 492264
rect 576509 493182 576567 493223
rect 576509 493148 576521 493182
rect 576555 493148 576567 493182
rect 576509 493114 576567 493148
rect 576509 493080 576521 493114
rect 576555 493080 576567 493114
rect 576509 493046 576567 493080
rect 576509 493012 576521 493046
rect 576555 493012 576567 493046
rect 576509 492978 576567 493012
rect 576509 492944 576521 492978
rect 576555 492944 576567 492978
rect 576509 492910 576567 492944
rect 576509 492876 576521 492910
rect 576555 492876 576567 492910
rect 576509 492842 576567 492876
rect 576509 492808 576521 492842
rect 576555 492808 576567 492842
rect 576509 492774 576567 492808
rect 576509 492740 576521 492774
rect 576555 492740 576567 492774
rect 576509 492706 576567 492740
rect 576509 492672 576521 492706
rect 576555 492672 576567 492706
rect 576509 492638 576567 492672
rect 576509 492604 576521 492638
rect 576555 492604 576567 492638
rect 576509 492570 576567 492604
rect 576509 492536 576521 492570
rect 576555 492536 576567 492570
rect 576509 492502 576567 492536
rect 576509 492468 576521 492502
rect 576555 492468 576567 492502
rect 576509 492434 576567 492468
rect 576509 492400 576521 492434
rect 576555 492400 576567 492434
rect 576509 492366 576567 492400
rect 576509 492332 576521 492366
rect 576555 492332 576567 492366
rect 576509 492298 576567 492332
rect 576509 492264 576521 492298
rect 576555 492264 576567 492298
rect 576509 492223 576567 492264
rect 576767 493182 576825 493223
rect 576767 493148 576779 493182
rect 576813 493148 576825 493182
rect 576767 493114 576825 493148
rect 576767 493080 576779 493114
rect 576813 493080 576825 493114
rect 576767 493046 576825 493080
rect 576767 493012 576779 493046
rect 576813 493012 576825 493046
rect 576767 492978 576825 493012
rect 576767 492944 576779 492978
rect 576813 492944 576825 492978
rect 576767 492910 576825 492944
rect 576767 492876 576779 492910
rect 576813 492876 576825 492910
rect 576767 492842 576825 492876
rect 576767 492808 576779 492842
rect 576813 492808 576825 492842
rect 576767 492774 576825 492808
rect 576767 492740 576779 492774
rect 576813 492740 576825 492774
rect 576767 492706 576825 492740
rect 576767 492672 576779 492706
rect 576813 492672 576825 492706
rect 576767 492638 576825 492672
rect 576767 492604 576779 492638
rect 576813 492604 576825 492638
rect 576767 492570 576825 492604
rect 576767 492536 576779 492570
rect 576813 492536 576825 492570
rect 576767 492502 576825 492536
rect 576767 492468 576779 492502
rect 576813 492468 576825 492502
rect 576767 492434 576825 492468
rect 576767 492400 576779 492434
rect 576813 492400 576825 492434
rect 576767 492366 576825 492400
rect 576767 492332 576779 492366
rect 576813 492332 576825 492366
rect 576767 492298 576825 492332
rect 576767 492264 576779 492298
rect 576813 492264 576825 492298
rect 576767 492223 576825 492264
rect 577025 493182 577083 493223
rect 577025 493148 577037 493182
rect 577071 493148 577083 493182
rect 577025 493114 577083 493148
rect 577025 493080 577037 493114
rect 577071 493080 577083 493114
rect 577025 493046 577083 493080
rect 577025 493012 577037 493046
rect 577071 493012 577083 493046
rect 577025 492978 577083 493012
rect 577025 492944 577037 492978
rect 577071 492944 577083 492978
rect 577025 492910 577083 492944
rect 577025 492876 577037 492910
rect 577071 492876 577083 492910
rect 577025 492842 577083 492876
rect 577025 492808 577037 492842
rect 577071 492808 577083 492842
rect 577025 492774 577083 492808
rect 577025 492740 577037 492774
rect 577071 492740 577083 492774
rect 577025 492706 577083 492740
rect 577025 492672 577037 492706
rect 577071 492672 577083 492706
rect 577025 492638 577083 492672
rect 577025 492604 577037 492638
rect 577071 492604 577083 492638
rect 577025 492570 577083 492604
rect 577025 492536 577037 492570
rect 577071 492536 577083 492570
rect 577025 492502 577083 492536
rect 577025 492468 577037 492502
rect 577071 492468 577083 492502
rect 577025 492434 577083 492468
rect 577025 492400 577037 492434
rect 577071 492400 577083 492434
rect 577025 492366 577083 492400
rect 577025 492332 577037 492366
rect 577071 492332 577083 492366
rect 577025 492298 577083 492332
rect 577025 492264 577037 492298
rect 577071 492264 577083 492298
rect 577025 492223 577083 492264
rect 577283 493182 577341 493223
rect 577283 493148 577295 493182
rect 577329 493148 577341 493182
rect 577283 493114 577341 493148
rect 577283 493080 577295 493114
rect 577329 493080 577341 493114
rect 577283 493046 577341 493080
rect 577283 493012 577295 493046
rect 577329 493012 577341 493046
rect 577283 492978 577341 493012
rect 577283 492944 577295 492978
rect 577329 492944 577341 492978
rect 577283 492910 577341 492944
rect 577283 492876 577295 492910
rect 577329 492876 577341 492910
rect 577283 492842 577341 492876
rect 577283 492808 577295 492842
rect 577329 492808 577341 492842
rect 577283 492774 577341 492808
rect 577283 492740 577295 492774
rect 577329 492740 577341 492774
rect 577283 492706 577341 492740
rect 577283 492672 577295 492706
rect 577329 492672 577341 492706
rect 577283 492638 577341 492672
rect 577283 492604 577295 492638
rect 577329 492604 577341 492638
rect 577283 492570 577341 492604
rect 577283 492536 577295 492570
rect 577329 492536 577341 492570
rect 577283 492502 577341 492536
rect 577283 492468 577295 492502
rect 577329 492468 577341 492502
rect 577283 492434 577341 492468
rect 577283 492400 577295 492434
rect 577329 492400 577341 492434
rect 577283 492366 577341 492400
rect 577283 492332 577295 492366
rect 577329 492332 577341 492366
rect 577283 492298 577341 492332
rect 577283 492264 577295 492298
rect 577329 492264 577341 492298
rect 577283 492223 577341 492264
rect 577541 493182 577599 493223
rect 577541 493148 577553 493182
rect 577587 493148 577599 493182
rect 577541 493114 577599 493148
rect 577541 493080 577553 493114
rect 577587 493080 577599 493114
rect 577541 493046 577599 493080
rect 577541 493012 577553 493046
rect 577587 493012 577599 493046
rect 577541 492978 577599 493012
rect 577541 492944 577553 492978
rect 577587 492944 577599 492978
rect 577541 492910 577599 492944
rect 577541 492876 577553 492910
rect 577587 492876 577599 492910
rect 577541 492842 577599 492876
rect 577541 492808 577553 492842
rect 577587 492808 577599 492842
rect 577541 492774 577599 492808
rect 577541 492740 577553 492774
rect 577587 492740 577599 492774
rect 577541 492706 577599 492740
rect 577541 492672 577553 492706
rect 577587 492672 577599 492706
rect 577541 492638 577599 492672
rect 577541 492604 577553 492638
rect 577587 492604 577599 492638
rect 577541 492570 577599 492604
rect 577541 492536 577553 492570
rect 577587 492536 577599 492570
rect 577541 492502 577599 492536
rect 577541 492468 577553 492502
rect 577587 492468 577599 492502
rect 577541 492434 577599 492468
rect 577541 492400 577553 492434
rect 577587 492400 577599 492434
rect 577541 492366 577599 492400
rect 577541 492332 577553 492366
rect 577587 492332 577599 492366
rect 577541 492298 577599 492332
rect 577541 492264 577553 492298
rect 577587 492264 577599 492298
rect 577541 492223 577599 492264
rect 577799 493182 577857 493223
rect 577799 493148 577811 493182
rect 577845 493148 577857 493182
rect 577799 493114 577857 493148
rect 577799 493080 577811 493114
rect 577845 493080 577857 493114
rect 577799 493046 577857 493080
rect 577799 493012 577811 493046
rect 577845 493012 577857 493046
rect 577799 492978 577857 493012
rect 577799 492944 577811 492978
rect 577845 492944 577857 492978
rect 577799 492910 577857 492944
rect 577799 492876 577811 492910
rect 577845 492876 577857 492910
rect 577799 492842 577857 492876
rect 577799 492808 577811 492842
rect 577845 492808 577857 492842
rect 577799 492774 577857 492808
rect 577799 492740 577811 492774
rect 577845 492740 577857 492774
rect 577799 492706 577857 492740
rect 577799 492672 577811 492706
rect 577845 492672 577857 492706
rect 577799 492638 577857 492672
rect 577799 492604 577811 492638
rect 577845 492604 577857 492638
rect 577799 492570 577857 492604
rect 577799 492536 577811 492570
rect 577845 492536 577857 492570
rect 577799 492502 577857 492536
rect 577799 492468 577811 492502
rect 577845 492468 577857 492502
rect 577799 492434 577857 492468
rect 577799 492400 577811 492434
rect 577845 492400 577857 492434
rect 577799 492366 577857 492400
rect 577799 492332 577811 492366
rect 577845 492332 577857 492366
rect 577799 492298 577857 492332
rect 577799 492264 577811 492298
rect 577845 492264 577857 492298
rect 577799 492223 577857 492264
rect 578057 493182 578115 493223
rect 578057 493148 578069 493182
rect 578103 493148 578115 493182
rect 578057 493114 578115 493148
rect 578057 493080 578069 493114
rect 578103 493080 578115 493114
rect 578057 493046 578115 493080
rect 578057 493012 578069 493046
rect 578103 493012 578115 493046
rect 578057 492978 578115 493012
rect 578057 492944 578069 492978
rect 578103 492944 578115 492978
rect 578057 492910 578115 492944
rect 578057 492876 578069 492910
rect 578103 492876 578115 492910
rect 578057 492842 578115 492876
rect 578057 492808 578069 492842
rect 578103 492808 578115 492842
rect 578057 492774 578115 492808
rect 578057 492740 578069 492774
rect 578103 492740 578115 492774
rect 578057 492706 578115 492740
rect 578057 492672 578069 492706
rect 578103 492672 578115 492706
rect 578057 492638 578115 492672
rect 578057 492604 578069 492638
rect 578103 492604 578115 492638
rect 578057 492570 578115 492604
rect 578057 492536 578069 492570
rect 578103 492536 578115 492570
rect 578057 492502 578115 492536
rect 578057 492468 578069 492502
rect 578103 492468 578115 492502
rect 578057 492434 578115 492468
rect 578057 492400 578069 492434
rect 578103 492400 578115 492434
rect 578057 492366 578115 492400
rect 578057 492332 578069 492366
rect 578103 492332 578115 492366
rect 578057 492298 578115 492332
rect 578057 492264 578069 492298
rect 578103 492264 578115 492298
rect 578057 492223 578115 492264
rect 578315 493182 578373 493223
rect 578315 493148 578327 493182
rect 578361 493148 578373 493182
rect 578315 493114 578373 493148
rect 578315 493080 578327 493114
rect 578361 493080 578373 493114
rect 578315 493046 578373 493080
rect 578315 493012 578327 493046
rect 578361 493012 578373 493046
rect 578315 492978 578373 493012
rect 578315 492944 578327 492978
rect 578361 492944 578373 492978
rect 578315 492910 578373 492944
rect 578315 492876 578327 492910
rect 578361 492876 578373 492910
rect 578315 492842 578373 492876
rect 578315 492808 578327 492842
rect 578361 492808 578373 492842
rect 578315 492774 578373 492808
rect 578315 492740 578327 492774
rect 578361 492740 578373 492774
rect 578315 492706 578373 492740
rect 578315 492672 578327 492706
rect 578361 492672 578373 492706
rect 578315 492638 578373 492672
rect 578315 492604 578327 492638
rect 578361 492604 578373 492638
rect 578315 492570 578373 492604
rect 578315 492536 578327 492570
rect 578361 492536 578373 492570
rect 578315 492502 578373 492536
rect 578315 492468 578327 492502
rect 578361 492468 578373 492502
rect 578315 492434 578373 492468
rect 578315 492400 578327 492434
rect 578361 492400 578373 492434
rect 578315 492366 578373 492400
rect 578315 492332 578327 492366
rect 578361 492332 578373 492366
rect 578315 492298 578373 492332
rect 578315 492264 578327 492298
rect 578361 492264 578373 492298
rect 578315 492223 578373 492264
rect 578573 493182 578631 493223
rect 578573 493148 578585 493182
rect 578619 493148 578631 493182
rect 578573 493114 578631 493148
rect 578573 493080 578585 493114
rect 578619 493080 578631 493114
rect 578573 493046 578631 493080
rect 578573 493012 578585 493046
rect 578619 493012 578631 493046
rect 578573 492978 578631 493012
rect 578573 492944 578585 492978
rect 578619 492944 578631 492978
rect 578573 492910 578631 492944
rect 578573 492876 578585 492910
rect 578619 492876 578631 492910
rect 578573 492842 578631 492876
rect 578573 492808 578585 492842
rect 578619 492808 578631 492842
rect 578573 492774 578631 492808
rect 578573 492740 578585 492774
rect 578619 492740 578631 492774
rect 578573 492706 578631 492740
rect 578573 492672 578585 492706
rect 578619 492672 578631 492706
rect 578573 492638 578631 492672
rect 578573 492604 578585 492638
rect 578619 492604 578631 492638
rect 578573 492570 578631 492604
rect 578573 492536 578585 492570
rect 578619 492536 578631 492570
rect 578573 492502 578631 492536
rect 578573 492468 578585 492502
rect 578619 492468 578631 492502
rect 578573 492434 578631 492468
rect 578573 492400 578585 492434
rect 578619 492400 578631 492434
rect 578573 492366 578631 492400
rect 578573 492332 578585 492366
rect 578619 492332 578631 492366
rect 578573 492298 578631 492332
rect 578573 492264 578585 492298
rect 578619 492264 578631 492298
rect 578573 492223 578631 492264
rect 578831 493182 578889 493223
rect 578831 493148 578843 493182
rect 578877 493148 578889 493182
rect 578831 493114 578889 493148
rect 578831 493080 578843 493114
rect 578877 493080 578889 493114
rect 578831 493046 578889 493080
rect 578831 493012 578843 493046
rect 578877 493012 578889 493046
rect 578831 492978 578889 493012
rect 578831 492944 578843 492978
rect 578877 492944 578889 492978
rect 578831 492910 578889 492944
rect 578831 492876 578843 492910
rect 578877 492876 578889 492910
rect 578831 492842 578889 492876
rect 578831 492808 578843 492842
rect 578877 492808 578889 492842
rect 578831 492774 578889 492808
rect 578831 492740 578843 492774
rect 578877 492740 578889 492774
rect 578831 492706 578889 492740
rect 578831 492672 578843 492706
rect 578877 492672 578889 492706
rect 578831 492638 578889 492672
rect 578831 492604 578843 492638
rect 578877 492604 578889 492638
rect 578831 492570 578889 492604
rect 578831 492536 578843 492570
rect 578877 492536 578889 492570
rect 578831 492502 578889 492536
rect 578831 492468 578843 492502
rect 578877 492468 578889 492502
rect 578831 492434 578889 492468
rect 578831 492400 578843 492434
rect 578877 492400 578889 492434
rect 578831 492366 578889 492400
rect 578831 492332 578843 492366
rect 578877 492332 578889 492366
rect 578831 492298 578889 492332
rect 578831 492264 578843 492298
rect 578877 492264 578889 492298
rect 578831 492223 578889 492264
rect 579089 493182 579147 493223
rect 579089 493148 579101 493182
rect 579135 493148 579147 493182
rect 579089 493114 579147 493148
rect 579089 493080 579101 493114
rect 579135 493080 579147 493114
rect 579089 493046 579147 493080
rect 579089 493012 579101 493046
rect 579135 493012 579147 493046
rect 579089 492978 579147 493012
rect 579089 492944 579101 492978
rect 579135 492944 579147 492978
rect 579089 492910 579147 492944
rect 579089 492876 579101 492910
rect 579135 492876 579147 492910
rect 579089 492842 579147 492876
rect 579089 492808 579101 492842
rect 579135 492808 579147 492842
rect 579089 492774 579147 492808
rect 579089 492740 579101 492774
rect 579135 492740 579147 492774
rect 579089 492706 579147 492740
rect 579089 492672 579101 492706
rect 579135 492672 579147 492706
rect 579089 492638 579147 492672
rect 579089 492604 579101 492638
rect 579135 492604 579147 492638
rect 579089 492570 579147 492604
rect 579089 492536 579101 492570
rect 579135 492536 579147 492570
rect 579089 492502 579147 492536
rect 579089 492468 579101 492502
rect 579135 492468 579147 492502
rect 579089 492434 579147 492468
rect 579089 492400 579101 492434
rect 579135 492400 579147 492434
rect 579089 492366 579147 492400
rect 579089 492332 579101 492366
rect 579135 492332 579147 492366
rect 579089 492298 579147 492332
rect 579089 492264 579101 492298
rect 579135 492264 579147 492298
rect 579089 492223 579147 492264
rect 579347 493182 579405 493223
rect 579347 493148 579359 493182
rect 579393 493148 579405 493182
rect 579347 493114 579405 493148
rect 579347 493080 579359 493114
rect 579393 493080 579405 493114
rect 579347 493046 579405 493080
rect 579347 493012 579359 493046
rect 579393 493012 579405 493046
rect 579347 492978 579405 493012
rect 579347 492944 579359 492978
rect 579393 492944 579405 492978
rect 579347 492910 579405 492944
rect 579347 492876 579359 492910
rect 579393 492876 579405 492910
rect 579347 492842 579405 492876
rect 579347 492808 579359 492842
rect 579393 492808 579405 492842
rect 579347 492774 579405 492808
rect 579347 492740 579359 492774
rect 579393 492740 579405 492774
rect 579347 492706 579405 492740
rect 579347 492672 579359 492706
rect 579393 492672 579405 492706
rect 579347 492638 579405 492672
rect 579347 492604 579359 492638
rect 579393 492604 579405 492638
rect 579347 492570 579405 492604
rect 579347 492536 579359 492570
rect 579393 492536 579405 492570
rect 579347 492502 579405 492536
rect 579347 492468 579359 492502
rect 579393 492468 579405 492502
rect 579347 492434 579405 492468
rect 579347 492400 579359 492434
rect 579393 492400 579405 492434
rect 579347 492366 579405 492400
rect 579347 492332 579359 492366
rect 579393 492332 579405 492366
rect 579347 492298 579405 492332
rect 579347 492264 579359 492298
rect 579393 492264 579405 492298
rect 579347 492223 579405 492264
rect 579605 493182 579663 493223
rect 579605 493148 579617 493182
rect 579651 493148 579663 493182
rect 579605 493114 579663 493148
rect 579605 493080 579617 493114
rect 579651 493080 579663 493114
rect 579605 493046 579663 493080
rect 579605 493012 579617 493046
rect 579651 493012 579663 493046
rect 579605 492978 579663 493012
rect 579605 492944 579617 492978
rect 579651 492944 579663 492978
rect 579605 492910 579663 492944
rect 579605 492876 579617 492910
rect 579651 492876 579663 492910
rect 579605 492842 579663 492876
rect 579605 492808 579617 492842
rect 579651 492808 579663 492842
rect 579605 492774 579663 492808
rect 579605 492740 579617 492774
rect 579651 492740 579663 492774
rect 579605 492706 579663 492740
rect 579605 492672 579617 492706
rect 579651 492672 579663 492706
rect 579605 492638 579663 492672
rect 579605 492604 579617 492638
rect 579651 492604 579663 492638
rect 579605 492570 579663 492604
rect 579605 492536 579617 492570
rect 579651 492536 579663 492570
rect 579605 492502 579663 492536
rect 579605 492468 579617 492502
rect 579651 492468 579663 492502
rect 579605 492434 579663 492468
rect 579605 492400 579617 492434
rect 579651 492400 579663 492434
rect 579605 492366 579663 492400
rect 579605 492332 579617 492366
rect 579651 492332 579663 492366
rect 579605 492298 579663 492332
rect 579605 492264 579617 492298
rect 579651 492264 579663 492298
rect 579605 492223 579663 492264
rect 579863 493182 579921 493223
rect 579863 493148 579875 493182
rect 579909 493148 579921 493182
rect 579863 493114 579921 493148
rect 579863 493080 579875 493114
rect 579909 493080 579921 493114
rect 579863 493046 579921 493080
rect 579863 493012 579875 493046
rect 579909 493012 579921 493046
rect 579863 492978 579921 493012
rect 579863 492944 579875 492978
rect 579909 492944 579921 492978
rect 579863 492910 579921 492944
rect 579863 492876 579875 492910
rect 579909 492876 579921 492910
rect 579863 492842 579921 492876
rect 579863 492808 579875 492842
rect 579909 492808 579921 492842
rect 579863 492774 579921 492808
rect 579863 492740 579875 492774
rect 579909 492740 579921 492774
rect 579863 492706 579921 492740
rect 579863 492672 579875 492706
rect 579909 492672 579921 492706
rect 579863 492638 579921 492672
rect 579863 492604 579875 492638
rect 579909 492604 579921 492638
rect 579863 492570 579921 492604
rect 579863 492536 579875 492570
rect 579909 492536 579921 492570
rect 579863 492502 579921 492536
rect 579863 492468 579875 492502
rect 579909 492468 579921 492502
rect 579863 492434 579921 492468
rect 579863 492400 579875 492434
rect 579909 492400 579921 492434
rect 579863 492366 579921 492400
rect 579863 492332 579875 492366
rect 579909 492332 579921 492366
rect 579863 492298 579921 492332
rect 579863 492264 579875 492298
rect 579909 492264 579921 492298
rect 579863 492223 579921 492264
rect 580121 493182 580179 493223
rect 580121 493148 580133 493182
rect 580167 493148 580179 493182
rect 580121 493114 580179 493148
rect 580121 493080 580133 493114
rect 580167 493080 580179 493114
rect 580121 493046 580179 493080
rect 580121 493012 580133 493046
rect 580167 493012 580179 493046
rect 580121 492978 580179 493012
rect 580121 492944 580133 492978
rect 580167 492944 580179 492978
rect 580121 492910 580179 492944
rect 580121 492876 580133 492910
rect 580167 492876 580179 492910
rect 580121 492842 580179 492876
rect 580121 492808 580133 492842
rect 580167 492808 580179 492842
rect 580121 492774 580179 492808
rect 580121 492740 580133 492774
rect 580167 492740 580179 492774
rect 580121 492706 580179 492740
rect 580121 492672 580133 492706
rect 580167 492672 580179 492706
rect 580121 492638 580179 492672
rect 580121 492604 580133 492638
rect 580167 492604 580179 492638
rect 580121 492570 580179 492604
rect 580121 492536 580133 492570
rect 580167 492536 580179 492570
rect 580121 492502 580179 492536
rect 580121 492468 580133 492502
rect 580167 492468 580179 492502
rect 580121 492434 580179 492468
rect 580121 492400 580133 492434
rect 580167 492400 580179 492434
rect 580121 492366 580179 492400
rect 580121 492332 580133 492366
rect 580167 492332 580179 492366
rect 580121 492298 580179 492332
rect 580121 492264 580133 492298
rect 580167 492264 580179 492298
rect 580121 492223 580179 492264
rect 580379 493182 580437 493223
rect 580379 493148 580391 493182
rect 580425 493148 580437 493182
rect 580379 493114 580437 493148
rect 580379 493080 580391 493114
rect 580425 493080 580437 493114
rect 580379 493046 580437 493080
rect 580379 493012 580391 493046
rect 580425 493012 580437 493046
rect 580379 492978 580437 493012
rect 580379 492944 580391 492978
rect 580425 492944 580437 492978
rect 580379 492910 580437 492944
rect 580379 492876 580391 492910
rect 580425 492876 580437 492910
rect 580379 492842 580437 492876
rect 580379 492808 580391 492842
rect 580425 492808 580437 492842
rect 580379 492774 580437 492808
rect 580379 492740 580391 492774
rect 580425 492740 580437 492774
rect 580379 492706 580437 492740
rect 580379 492672 580391 492706
rect 580425 492672 580437 492706
rect 580379 492638 580437 492672
rect 580379 492604 580391 492638
rect 580425 492604 580437 492638
rect 580379 492570 580437 492604
rect 580379 492536 580391 492570
rect 580425 492536 580437 492570
rect 580379 492502 580437 492536
rect 580379 492468 580391 492502
rect 580425 492468 580437 492502
rect 580379 492434 580437 492468
rect 580379 492400 580391 492434
rect 580425 492400 580437 492434
rect 580379 492366 580437 492400
rect 580379 492332 580391 492366
rect 580425 492332 580437 492366
rect 580379 492298 580437 492332
rect 580379 492264 580391 492298
rect 580425 492264 580437 492298
rect 580379 492223 580437 492264
rect 574693 358878 574751 358919
rect 574693 358844 574705 358878
rect 574739 358844 574751 358878
rect 574693 358810 574751 358844
rect 574693 358776 574705 358810
rect 574739 358776 574751 358810
rect 574693 358742 574751 358776
rect 574693 358708 574705 358742
rect 574739 358708 574751 358742
rect 574693 358674 574751 358708
rect 574693 358640 574705 358674
rect 574739 358640 574751 358674
rect 574693 358606 574751 358640
rect 574693 358572 574705 358606
rect 574739 358572 574751 358606
rect 574693 358538 574751 358572
rect 574693 358504 574705 358538
rect 574739 358504 574751 358538
rect 574693 358470 574751 358504
rect 574693 358436 574705 358470
rect 574739 358436 574751 358470
rect 574693 358402 574751 358436
rect 574693 358368 574705 358402
rect 574739 358368 574751 358402
rect 574693 358334 574751 358368
rect 574693 358300 574705 358334
rect 574739 358300 574751 358334
rect 574693 358266 574751 358300
rect 574693 358232 574705 358266
rect 574739 358232 574751 358266
rect 574693 358198 574751 358232
rect 574693 358164 574705 358198
rect 574739 358164 574751 358198
rect 574693 358130 574751 358164
rect 574693 358096 574705 358130
rect 574739 358096 574751 358130
rect 574693 358062 574751 358096
rect 574693 358028 574705 358062
rect 574739 358028 574751 358062
rect 574693 357994 574751 358028
rect 574693 357960 574705 357994
rect 574739 357960 574751 357994
rect 574693 357919 574751 357960
rect 574951 358878 575009 358919
rect 574951 358844 574963 358878
rect 574997 358844 575009 358878
rect 574951 358810 575009 358844
rect 574951 358776 574963 358810
rect 574997 358776 575009 358810
rect 574951 358742 575009 358776
rect 574951 358708 574963 358742
rect 574997 358708 575009 358742
rect 574951 358674 575009 358708
rect 574951 358640 574963 358674
rect 574997 358640 575009 358674
rect 574951 358606 575009 358640
rect 574951 358572 574963 358606
rect 574997 358572 575009 358606
rect 574951 358538 575009 358572
rect 574951 358504 574963 358538
rect 574997 358504 575009 358538
rect 574951 358470 575009 358504
rect 574951 358436 574963 358470
rect 574997 358436 575009 358470
rect 574951 358402 575009 358436
rect 574951 358368 574963 358402
rect 574997 358368 575009 358402
rect 574951 358334 575009 358368
rect 574951 358300 574963 358334
rect 574997 358300 575009 358334
rect 574951 358266 575009 358300
rect 574951 358232 574963 358266
rect 574997 358232 575009 358266
rect 574951 358198 575009 358232
rect 574951 358164 574963 358198
rect 574997 358164 575009 358198
rect 574951 358130 575009 358164
rect 574951 358096 574963 358130
rect 574997 358096 575009 358130
rect 574951 358062 575009 358096
rect 574951 358028 574963 358062
rect 574997 358028 575009 358062
rect 574951 357994 575009 358028
rect 574951 357960 574963 357994
rect 574997 357960 575009 357994
rect 574951 357919 575009 357960
rect 575209 358878 575267 358919
rect 575209 358844 575221 358878
rect 575255 358844 575267 358878
rect 575209 358810 575267 358844
rect 575209 358776 575221 358810
rect 575255 358776 575267 358810
rect 575209 358742 575267 358776
rect 575209 358708 575221 358742
rect 575255 358708 575267 358742
rect 575209 358674 575267 358708
rect 575209 358640 575221 358674
rect 575255 358640 575267 358674
rect 575209 358606 575267 358640
rect 575209 358572 575221 358606
rect 575255 358572 575267 358606
rect 575209 358538 575267 358572
rect 575209 358504 575221 358538
rect 575255 358504 575267 358538
rect 575209 358470 575267 358504
rect 575209 358436 575221 358470
rect 575255 358436 575267 358470
rect 575209 358402 575267 358436
rect 575209 358368 575221 358402
rect 575255 358368 575267 358402
rect 575209 358334 575267 358368
rect 575209 358300 575221 358334
rect 575255 358300 575267 358334
rect 575209 358266 575267 358300
rect 575209 358232 575221 358266
rect 575255 358232 575267 358266
rect 575209 358198 575267 358232
rect 575209 358164 575221 358198
rect 575255 358164 575267 358198
rect 575209 358130 575267 358164
rect 575209 358096 575221 358130
rect 575255 358096 575267 358130
rect 575209 358062 575267 358096
rect 575209 358028 575221 358062
rect 575255 358028 575267 358062
rect 575209 357994 575267 358028
rect 575209 357960 575221 357994
rect 575255 357960 575267 357994
rect 575209 357919 575267 357960
rect 575467 358878 575525 358919
rect 575467 358844 575479 358878
rect 575513 358844 575525 358878
rect 575467 358810 575525 358844
rect 575467 358776 575479 358810
rect 575513 358776 575525 358810
rect 575467 358742 575525 358776
rect 575467 358708 575479 358742
rect 575513 358708 575525 358742
rect 575467 358674 575525 358708
rect 575467 358640 575479 358674
rect 575513 358640 575525 358674
rect 575467 358606 575525 358640
rect 575467 358572 575479 358606
rect 575513 358572 575525 358606
rect 575467 358538 575525 358572
rect 575467 358504 575479 358538
rect 575513 358504 575525 358538
rect 575467 358470 575525 358504
rect 575467 358436 575479 358470
rect 575513 358436 575525 358470
rect 575467 358402 575525 358436
rect 575467 358368 575479 358402
rect 575513 358368 575525 358402
rect 575467 358334 575525 358368
rect 575467 358300 575479 358334
rect 575513 358300 575525 358334
rect 575467 358266 575525 358300
rect 575467 358232 575479 358266
rect 575513 358232 575525 358266
rect 575467 358198 575525 358232
rect 575467 358164 575479 358198
rect 575513 358164 575525 358198
rect 575467 358130 575525 358164
rect 575467 358096 575479 358130
rect 575513 358096 575525 358130
rect 575467 358062 575525 358096
rect 575467 358028 575479 358062
rect 575513 358028 575525 358062
rect 575467 357994 575525 358028
rect 575467 357960 575479 357994
rect 575513 357960 575525 357994
rect 575467 357919 575525 357960
rect 575725 358878 575783 358919
rect 575725 358844 575737 358878
rect 575771 358844 575783 358878
rect 575725 358810 575783 358844
rect 575725 358776 575737 358810
rect 575771 358776 575783 358810
rect 575725 358742 575783 358776
rect 575725 358708 575737 358742
rect 575771 358708 575783 358742
rect 575725 358674 575783 358708
rect 575725 358640 575737 358674
rect 575771 358640 575783 358674
rect 575725 358606 575783 358640
rect 575725 358572 575737 358606
rect 575771 358572 575783 358606
rect 575725 358538 575783 358572
rect 575725 358504 575737 358538
rect 575771 358504 575783 358538
rect 575725 358470 575783 358504
rect 575725 358436 575737 358470
rect 575771 358436 575783 358470
rect 575725 358402 575783 358436
rect 575725 358368 575737 358402
rect 575771 358368 575783 358402
rect 575725 358334 575783 358368
rect 575725 358300 575737 358334
rect 575771 358300 575783 358334
rect 575725 358266 575783 358300
rect 575725 358232 575737 358266
rect 575771 358232 575783 358266
rect 575725 358198 575783 358232
rect 575725 358164 575737 358198
rect 575771 358164 575783 358198
rect 575725 358130 575783 358164
rect 575725 358096 575737 358130
rect 575771 358096 575783 358130
rect 575725 358062 575783 358096
rect 575725 358028 575737 358062
rect 575771 358028 575783 358062
rect 575725 357994 575783 358028
rect 575725 357960 575737 357994
rect 575771 357960 575783 357994
rect 575725 357919 575783 357960
rect 575983 358878 576041 358919
rect 575983 358844 575995 358878
rect 576029 358844 576041 358878
rect 575983 358810 576041 358844
rect 575983 358776 575995 358810
rect 576029 358776 576041 358810
rect 575983 358742 576041 358776
rect 575983 358708 575995 358742
rect 576029 358708 576041 358742
rect 575983 358674 576041 358708
rect 575983 358640 575995 358674
rect 576029 358640 576041 358674
rect 575983 358606 576041 358640
rect 575983 358572 575995 358606
rect 576029 358572 576041 358606
rect 575983 358538 576041 358572
rect 575983 358504 575995 358538
rect 576029 358504 576041 358538
rect 575983 358470 576041 358504
rect 575983 358436 575995 358470
rect 576029 358436 576041 358470
rect 575983 358402 576041 358436
rect 575983 358368 575995 358402
rect 576029 358368 576041 358402
rect 575983 358334 576041 358368
rect 575983 358300 575995 358334
rect 576029 358300 576041 358334
rect 575983 358266 576041 358300
rect 575983 358232 575995 358266
rect 576029 358232 576041 358266
rect 575983 358198 576041 358232
rect 575983 358164 575995 358198
rect 576029 358164 576041 358198
rect 575983 358130 576041 358164
rect 575983 358096 575995 358130
rect 576029 358096 576041 358130
rect 575983 358062 576041 358096
rect 575983 358028 575995 358062
rect 576029 358028 576041 358062
rect 575983 357994 576041 358028
rect 575983 357960 575995 357994
rect 576029 357960 576041 357994
rect 575983 357919 576041 357960
rect 576241 358878 576299 358919
rect 576241 358844 576253 358878
rect 576287 358844 576299 358878
rect 576241 358810 576299 358844
rect 576241 358776 576253 358810
rect 576287 358776 576299 358810
rect 576241 358742 576299 358776
rect 576241 358708 576253 358742
rect 576287 358708 576299 358742
rect 576241 358674 576299 358708
rect 576241 358640 576253 358674
rect 576287 358640 576299 358674
rect 576241 358606 576299 358640
rect 576241 358572 576253 358606
rect 576287 358572 576299 358606
rect 576241 358538 576299 358572
rect 576241 358504 576253 358538
rect 576287 358504 576299 358538
rect 576241 358470 576299 358504
rect 576241 358436 576253 358470
rect 576287 358436 576299 358470
rect 576241 358402 576299 358436
rect 576241 358368 576253 358402
rect 576287 358368 576299 358402
rect 576241 358334 576299 358368
rect 576241 358300 576253 358334
rect 576287 358300 576299 358334
rect 576241 358266 576299 358300
rect 576241 358232 576253 358266
rect 576287 358232 576299 358266
rect 576241 358198 576299 358232
rect 576241 358164 576253 358198
rect 576287 358164 576299 358198
rect 576241 358130 576299 358164
rect 576241 358096 576253 358130
rect 576287 358096 576299 358130
rect 576241 358062 576299 358096
rect 576241 358028 576253 358062
rect 576287 358028 576299 358062
rect 576241 357994 576299 358028
rect 576241 357960 576253 357994
rect 576287 357960 576299 357994
rect 576241 357919 576299 357960
rect 576499 358878 576557 358919
rect 576499 358844 576511 358878
rect 576545 358844 576557 358878
rect 576499 358810 576557 358844
rect 576499 358776 576511 358810
rect 576545 358776 576557 358810
rect 576499 358742 576557 358776
rect 576499 358708 576511 358742
rect 576545 358708 576557 358742
rect 576499 358674 576557 358708
rect 576499 358640 576511 358674
rect 576545 358640 576557 358674
rect 576499 358606 576557 358640
rect 576499 358572 576511 358606
rect 576545 358572 576557 358606
rect 576499 358538 576557 358572
rect 576499 358504 576511 358538
rect 576545 358504 576557 358538
rect 576499 358470 576557 358504
rect 576499 358436 576511 358470
rect 576545 358436 576557 358470
rect 576499 358402 576557 358436
rect 576499 358368 576511 358402
rect 576545 358368 576557 358402
rect 576499 358334 576557 358368
rect 576499 358300 576511 358334
rect 576545 358300 576557 358334
rect 576499 358266 576557 358300
rect 576499 358232 576511 358266
rect 576545 358232 576557 358266
rect 576499 358198 576557 358232
rect 576499 358164 576511 358198
rect 576545 358164 576557 358198
rect 576499 358130 576557 358164
rect 576499 358096 576511 358130
rect 576545 358096 576557 358130
rect 576499 358062 576557 358096
rect 576499 358028 576511 358062
rect 576545 358028 576557 358062
rect 576499 357994 576557 358028
rect 576499 357960 576511 357994
rect 576545 357960 576557 357994
rect 576499 357919 576557 357960
rect 576757 358878 576815 358919
rect 576757 358844 576769 358878
rect 576803 358844 576815 358878
rect 576757 358810 576815 358844
rect 576757 358776 576769 358810
rect 576803 358776 576815 358810
rect 576757 358742 576815 358776
rect 576757 358708 576769 358742
rect 576803 358708 576815 358742
rect 576757 358674 576815 358708
rect 576757 358640 576769 358674
rect 576803 358640 576815 358674
rect 576757 358606 576815 358640
rect 576757 358572 576769 358606
rect 576803 358572 576815 358606
rect 576757 358538 576815 358572
rect 576757 358504 576769 358538
rect 576803 358504 576815 358538
rect 576757 358470 576815 358504
rect 576757 358436 576769 358470
rect 576803 358436 576815 358470
rect 576757 358402 576815 358436
rect 576757 358368 576769 358402
rect 576803 358368 576815 358402
rect 576757 358334 576815 358368
rect 576757 358300 576769 358334
rect 576803 358300 576815 358334
rect 576757 358266 576815 358300
rect 576757 358232 576769 358266
rect 576803 358232 576815 358266
rect 576757 358198 576815 358232
rect 576757 358164 576769 358198
rect 576803 358164 576815 358198
rect 576757 358130 576815 358164
rect 576757 358096 576769 358130
rect 576803 358096 576815 358130
rect 576757 358062 576815 358096
rect 576757 358028 576769 358062
rect 576803 358028 576815 358062
rect 576757 357994 576815 358028
rect 576757 357960 576769 357994
rect 576803 357960 576815 357994
rect 576757 357919 576815 357960
rect 577015 358878 577073 358919
rect 577015 358844 577027 358878
rect 577061 358844 577073 358878
rect 577015 358810 577073 358844
rect 577015 358776 577027 358810
rect 577061 358776 577073 358810
rect 577015 358742 577073 358776
rect 577015 358708 577027 358742
rect 577061 358708 577073 358742
rect 577015 358674 577073 358708
rect 577015 358640 577027 358674
rect 577061 358640 577073 358674
rect 577015 358606 577073 358640
rect 577015 358572 577027 358606
rect 577061 358572 577073 358606
rect 577015 358538 577073 358572
rect 577015 358504 577027 358538
rect 577061 358504 577073 358538
rect 577015 358470 577073 358504
rect 577015 358436 577027 358470
rect 577061 358436 577073 358470
rect 577015 358402 577073 358436
rect 577015 358368 577027 358402
rect 577061 358368 577073 358402
rect 577015 358334 577073 358368
rect 577015 358300 577027 358334
rect 577061 358300 577073 358334
rect 577015 358266 577073 358300
rect 577015 358232 577027 358266
rect 577061 358232 577073 358266
rect 577015 358198 577073 358232
rect 577015 358164 577027 358198
rect 577061 358164 577073 358198
rect 577015 358130 577073 358164
rect 577015 358096 577027 358130
rect 577061 358096 577073 358130
rect 577015 358062 577073 358096
rect 577015 358028 577027 358062
rect 577061 358028 577073 358062
rect 577015 357994 577073 358028
rect 577015 357960 577027 357994
rect 577061 357960 577073 357994
rect 577015 357919 577073 357960
rect 577273 358878 577331 358919
rect 577273 358844 577285 358878
rect 577319 358844 577331 358878
rect 577273 358810 577331 358844
rect 577273 358776 577285 358810
rect 577319 358776 577331 358810
rect 577273 358742 577331 358776
rect 577273 358708 577285 358742
rect 577319 358708 577331 358742
rect 577273 358674 577331 358708
rect 577273 358640 577285 358674
rect 577319 358640 577331 358674
rect 577273 358606 577331 358640
rect 577273 358572 577285 358606
rect 577319 358572 577331 358606
rect 577273 358538 577331 358572
rect 577273 358504 577285 358538
rect 577319 358504 577331 358538
rect 577273 358470 577331 358504
rect 577273 358436 577285 358470
rect 577319 358436 577331 358470
rect 577273 358402 577331 358436
rect 577273 358368 577285 358402
rect 577319 358368 577331 358402
rect 577273 358334 577331 358368
rect 577273 358300 577285 358334
rect 577319 358300 577331 358334
rect 577273 358266 577331 358300
rect 577273 358232 577285 358266
rect 577319 358232 577331 358266
rect 577273 358198 577331 358232
rect 577273 358164 577285 358198
rect 577319 358164 577331 358198
rect 577273 358130 577331 358164
rect 577273 358096 577285 358130
rect 577319 358096 577331 358130
rect 577273 358062 577331 358096
rect 577273 358028 577285 358062
rect 577319 358028 577331 358062
rect 577273 357994 577331 358028
rect 577273 357960 577285 357994
rect 577319 357960 577331 357994
rect 577273 357919 577331 357960
rect 577531 358878 577589 358919
rect 577531 358844 577543 358878
rect 577577 358844 577589 358878
rect 577531 358810 577589 358844
rect 577531 358776 577543 358810
rect 577577 358776 577589 358810
rect 577531 358742 577589 358776
rect 577531 358708 577543 358742
rect 577577 358708 577589 358742
rect 577531 358674 577589 358708
rect 577531 358640 577543 358674
rect 577577 358640 577589 358674
rect 577531 358606 577589 358640
rect 577531 358572 577543 358606
rect 577577 358572 577589 358606
rect 577531 358538 577589 358572
rect 577531 358504 577543 358538
rect 577577 358504 577589 358538
rect 577531 358470 577589 358504
rect 577531 358436 577543 358470
rect 577577 358436 577589 358470
rect 577531 358402 577589 358436
rect 577531 358368 577543 358402
rect 577577 358368 577589 358402
rect 577531 358334 577589 358368
rect 577531 358300 577543 358334
rect 577577 358300 577589 358334
rect 577531 358266 577589 358300
rect 577531 358232 577543 358266
rect 577577 358232 577589 358266
rect 577531 358198 577589 358232
rect 577531 358164 577543 358198
rect 577577 358164 577589 358198
rect 577531 358130 577589 358164
rect 577531 358096 577543 358130
rect 577577 358096 577589 358130
rect 577531 358062 577589 358096
rect 577531 358028 577543 358062
rect 577577 358028 577589 358062
rect 577531 357994 577589 358028
rect 577531 357960 577543 357994
rect 577577 357960 577589 357994
rect 577531 357919 577589 357960
rect 577789 358878 577847 358919
rect 577789 358844 577801 358878
rect 577835 358844 577847 358878
rect 577789 358810 577847 358844
rect 577789 358776 577801 358810
rect 577835 358776 577847 358810
rect 577789 358742 577847 358776
rect 577789 358708 577801 358742
rect 577835 358708 577847 358742
rect 577789 358674 577847 358708
rect 577789 358640 577801 358674
rect 577835 358640 577847 358674
rect 577789 358606 577847 358640
rect 577789 358572 577801 358606
rect 577835 358572 577847 358606
rect 577789 358538 577847 358572
rect 577789 358504 577801 358538
rect 577835 358504 577847 358538
rect 577789 358470 577847 358504
rect 577789 358436 577801 358470
rect 577835 358436 577847 358470
rect 577789 358402 577847 358436
rect 577789 358368 577801 358402
rect 577835 358368 577847 358402
rect 577789 358334 577847 358368
rect 577789 358300 577801 358334
rect 577835 358300 577847 358334
rect 577789 358266 577847 358300
rect 577789 358232 577801 358266
rect 577835 358232 577847 358266
rect 577789 358198 577847 358232
rect 577789 358164 577801 358198
rect 577835 358164 577847 358198
rect 577789 358130 577847 358164
rect 577789 358096 577801 358130
rect 577835 358096 577847 358130
rect 577789 358062 577847 358096
rect 577789 358028 577801 358062
rect 577835 358028 577847 358062
rect 577789 357994 577847 358028
rect 577789 357960 577801 357994
rect 577835 357960 577847 357994
rect 577789 357919 577847 357960
rect 578047 358878 578105 358919
rect 578047 358844 578059 358878
rect 578093 358844 578105 358878
rect 578047 358810 578105 358844
rect 578047 358776 578059 358810
rect 578093 358776 578105 358810
rect 578047 358742 578105 358776
rect 578047 358708 578059 358742
rect 578093 358708 578105 358742
rect 578047 358674 578105 358708
rect 578047 358640 578059 358674
rect 578093 358640 578105 358674
rect 578047 358606 578105 358640
rect 578047 358572 578059 358606
rect 578093 358572 578105 358606
rect 578047 358538 578105 358572
rect 578047 358504 578059 358538
rect 578093 358504 578105 358538
rect 578047 358470 578105 358504
rect 578047 358436 578059 358470
rect 578093 358436 578105 358470
rect 578047 358402 578105 358436
rect 578047 358368 578059 358402
rect 578093 358368 578105 358402
rect 578047 358334 578105 358368
rect 578047 358300 578059 358334
rect 578093 358300 578105 358334
rect 578047 358266 578105 358300
rect 578047 358232 578059 358266
rect 578093 358232 578105 358266
rect 578047 358198 578105 358232
rect 578047 358164 578059 358198
rect 578093 358164 578105 358198
rect 578047 358130 578105 358164
rect 578047 358096 578059 358130
rect 578093 358096 578105 358130
rect 578047 358062 578105 358096
rect 578047 358028 578059 358062
rect 578093 358028 578105 358062
rect 578047 357994 578105 358028
rect 578047 357960 578059 357994
rect 578093 357960 578105 357994
rect 578047 357919 578105 357960
rect 578305 358878 578363 358919
rect 578305 358844 578317 358878
rect 578351 358844 578363 358878
rect 578305 358810 578363 358844
rect 578305 358776 578317 358810
rect 578351 358776 578363 358810
rect 578305 358742 578363 358776
rect 578305 358708 578317 358742
rect 578351 358708 578363 358742
rect 578305 358674 578363 358708
rect 578305 358640 578317 358674
rect 578351 358640 578363 358674
rect 578305 358606 578363 358640
rect 578305 358572 578317 358606
rect 578351 358572 578363 358606
rect 578305 358538 578363 358572
rect 578305 358504 578317 358538
rect 578351 358504 578363 358538
rect 578305 358470 578363 358504
rect 578305 358436 578317 358470
rect 578351 358436 578363 358470
rect 578305 358402 578363 358436
rect 578305 358368 578317 358402
rect 578351 358368 578363 358402
rect 578305 358334 578363 358368
rect 578305 358300 578317 358334
rect 578351 358300 578363 358334
rect 578305 358266 578363 358300
rect 578305 358232 578317 358266
rect 578351 358232 578363 358266
rect 578305 358198 578363 358232
rect 578305 358164 578317 358198
rect 578351 358164 578363 358198
rect 578305 358130 578363 358164
rect 578305 358096 578317 358130
rect 578351 358096 578363 358130
rect 578305 358062 578363 358096
rect 578305 358028 578317 358062
rect 578351 358028 578363 358062
rect 578305 357994 578363 358028
rect 578305 357960 578317 357994
rect 578351 357960 578363 357994
rect 578305 357919 578363 357960
rect 578563 358878 578621 358919
rect 578563 358844 578575 358878
rect 578609 358844 578621 358878
rect 578563 358810 578621 358844
rect 578563 358776 578575 358810
rect 578609 358776 578621 358810
rect 578563 358742 578621 358776
rect 578563 358708 578575 358742
rect 578609 358708 578621 358742
rect 578563 358674 578621 358708
rect 578563 358640 578575 358674
rect 578609 358640 578621 358674
rect 578563 358606 578621 358640
rect 578563 358572 578575 358606
rect 578609 358572 578621 358606
rect 578563 358538 578621 358572
rect 578563 358504 578575 358538
rect 578609 358504 578621 358538
rect 578563 358470 578621 358504
rect 578563 358436 578575 358470
rect 578609 358436 578621 358470
rect 578563 358402 578621 358436
rect 578563 358368 578575 358402
rect 578609 358368 578621 358402
rect 578563 358334 578621 358368
rect 578563 358300 578575 358334
rect 578609 358300 578621 358334
rect 578563 358266 578621 358300
rect 578563 358232 578575 358266
rect 578609 358232 578621 358266
rect 578563 358198 578621 358232
rect 578563 358164 578575 358198
rect 578609 358164 578621 358198
rect 578563 358130 578621 358164
rect 578563 358096 578575 358130
rect 578609 358096 578621 358130
rect 578563 358062 578621 358096
rect 578563 358028 578575 358062
rect 578609 358028 578621 358062
rect 578563 357994 578621 358028
rect 578563 357960 578575 357994
rect 578609 357960 578621 357994
rect 578563 357919 578621 357960
rect 578821 358878 578879 358919
rect 578821 358844 578833 358878
rect 578867 358844 578879 358878
rect 578821 358810 578879 358844
rect 578821 358776 578833 358810
rect 578867 358776 578879 358810
rect 578821 358742 578879 358776
rect 578821 358708 578833 358742
rect 578867 358708 578879 358742
rect 578821 358674 578879 358708
rect 578821 358640 578833 358674
rect 578867 358640 578879 358674
rect 578821 358606 578879 358640
rect 578821 358572 578833 358606
rect 578867 358572 578879 358606
rect 578821 358538 578879 358572
rect 578821 358504 578833 358538
rect 578867 358504 578879 358538
rect 578821 358470 578879 358504
rect 578821 358436 578833 358470
rect 578867 358436 578879 358470
rect 578821 358402 578879 358436
rect 578821 358368 578833 358402
rect 578867 358368 578879 358402
rect 578821 358334 578879 358368
rect 578821 358300 578833 358334
rect 578867 358300 578879 358334
rect 578821 358266 578879 358300
rect 578821 358232 578833 358266
rect 578867 358232 578879 358266
rect 578821 358198 578879 358232
rect 578821 358164 578833 358198
rect 578867 358164 578879 358198
rect 578821 358130 578879 358164
rect 578821 358096 578833 358130
rect 578867 358096 578879 358130
rect 578821 358062 578879 358096
rect 578821 358028 578833 358062
rect 578867 358028 578879 358062
rect 578821 357994 578879 358028
rect 578821 357960 578833 357994
rect 578867 357960 578879 357994
rect 578821 357919 578879 357960
rect 579079 358878 579137 358919
rect 579079 358844 579091 358878
rect 579125 358844 579137 358878
rect 579079 358810 579137 358844
rect 579079 358776 579091 358810
rect 579125 358776 579137 358810
rect 579079 358742 579137 358776
rect 579079 358708 579091 358742
rect 579125 358708 579137 358742
rect 579079 358674 579137 358708
rect 579079 358640 579091 358674
rect 579125 358640 579137 358674
rect 579079 358606 579137 358640
rect 579079 358572 579091 358606
rect 579125 358572 579137 358606
rect 579079 358538 579137 358572
rect 579079 358504 579091 358538
rect 579125 358504 579137 358538
rect 579079 358470 579137 358504
rect 579079 358436 579091 358470
rect 579125 358436 579137 358470
rect 579079 358402 579137 358436
rect 579079 358368 579091 358402
rect 579125 358368 579137 358402
rect 579079 358334 579137 358368
rect 579079 358300 579091 358334
rect 579125 358300 579137 358334
rect 579079 358266 579137 358300
rect 579079 358232 579091 358266
rect 579125 358232 579137 358266
rect 579079 358198 579137 358232
rect 579079 358164 579091 358198
rect 579125 358164 579137 358198
rect 579079 358130 579137 358164
rect 579079 358096 579091 358130
rect 579125 358096 579137 358130
rect 579079 358062 579137 358096
rect 579079 358028 579091 358062
rect 579125 358028 579137 358062
rect 579079 357994 579137 358028
rect 579079 357960 579091 357994
rect 579125 357960 579137 357994
rect 579079 357919 579137 357960
rect 579337 358878 579395 358919
rect 579337 358844 579349 358878
rect 579383 358844 579395 358878
rect 579337 358810 579395 358844
rect 579337 358776 579349 358810
rect 579383 358776 579395 358810
rect 579337 358742 579395 358776
rect 579337 358708 579349 358742
rect 579383 358708 579395 358742
rect 579337 358674 579395 358708
rect 579337 358640 579349 358674
rect 579383 358640 579395 358674
rect 579337 358606 579395 358640
rect 579337 358572 579349 358606
rect 579383 358572 579395 358606
rect 579337 358538 579395 358572
rect 579337 358504 579349 358538
rect 579383 358504 579395 358538
rect 579337 358470 579395 358504
rect 579337 358436 579349 358470
rect 579383 358436 579395 358470
rect 579337 358402 579395 358436
rect 579337 358368 579349 358402
rect 579383 358368 579395 358402
rect 579337 358334 579395 358368
rect 579337 358300 579349 358334
rect 579383 358300 579395 358334
rect 579337 358266 579395 358300
rect 579337 358232 579349 358266
rect 579383 358232 579395 358266
rect 579337 358198 579395 358232
rect 579337 358164 579349 358198
rect 579383 358164 579395 358198
rect 579337 358130 579395 358164
rect 579337 358096 579349 358130
rect 579383 358096 579395 358130
rect 579337 358062 579395 358096
rect 579337 358028 579349 358062
rect 579383 358028 579395 358062
rect 579337 357994 579395 358028
rect 579337 357960 579349 357994
rect 579383 357960 579395 357994
rect 579337 357919 579395 357960
rect 579595 358878 579653 358919
rect 579595 358844 579607 358878
rect 579641 358844 579653 358878
rect 579595 358810 579653 358844
rect 579595 358776 579607 358810
rect 579641 358776 579653 358810
rect 579595 358742 579653 358776
rect 579595 358708 579607 358742
rect 579641 358708 579653 358742
rect 579595 358674 579653 358708
rect 579595 358640 579607 358674
rect 579641 358640 579653 358674
rect 579595 358606 579653 358640
rect 579595 358572 579607 358606
rect 579641 358572 579653 358606
rect 579595 358538 579653 358572
rect 579595 358504 579607 358538
rect 579641 358504 579653 358538
rect 579595 358470 579653 358504
rect 579595 358436 579607 358470
rect 579641 358436 579653 358470
rect 579595 358402 579653 358436
rect 579595 358368 579607 358402
rect 579641 358368 579653 358402
rect 579595 358334 579653 358368
rect 579595 358300 579607 358334
rect 579641 358300 579653 358334
rect 579595 358266 579653 358300
rect 579595 358232 579607 358266
rect 579641 358232 579653 358266
rect 579595 358198 579653 358232
rect 579595 358164 579607 358198
rect 579641 358164 579653 358198
rect 579595 358130 579653 358164
rect 579595 358096 579607 358130
rect 579641 358096 579653 358130
rect 579595 358062 579653 358096
rect 579595 358028 579607 358062
rect 579641 358028 579653 358062
rect 579595 357994 579653 358028
rect 579595 357960 579607 357994
rect 579641 357960 579653 357994
rect 579595 357919 579653 357960
rect 579853 358878 579911 358919
rect 579853 358844 579865 358878
rect 579899 358844 579911 358878
rect 579853 358810 579911 358844
rect 579853 358776 579865 358810
rect 579899 358776 579911 358810
rect 579853 358742 579911 358776
rect 579853 358708 579865 358742
rect 579899 358708 579911 358742
rect 579853 358674 579911 358708
rect 579853 358640 579865 358674
rect 579899 358640 579911 358674
rect 579853 358606 579911 358640
rect 579853 358572 579865 358606
rect 579899 358572 579911 358606
rect 579853 358538 579911 358572
rect 579853 358504 579865 358538
rect 579899 358504 579911 358538
rect 579853 358470 579911 358504
rect 579853 358436 579865 358470
rect 579899 358436 579911 358470
rect 579853 358402 579911 358436
rect 579853 358368 579865 358402
rect 579899 358368 579911 358402
rect 579853 358334 579911 358368
rect 579853 358300 579865 358334
rect 579899 358300 579911 358334
rect 579853 358266 579911 358300
rect 579853 358232 579865 358266
rect 579899 358232 579911 358266
rect 579853 358198 579911 358232
rect 579853 358164 579865 358198
rect 579899 358164 579911 358198
rect 579853 358130 579911 358164
rect 579853 358096 579865 358130
rect 579899 358096 579911 358130
rect 579853 358062 579911 358096
rect 579853 358028 579865 358062
rect 579899 358028 579911 358062
rect 579853 357994 579911 358028
rect 579853 357960 579865 357994
rect 579899 357960 579911 357994
rect 579853 357919 579911 357960
rect 575141 312710 575199 312751
rect 575141 312676 575153 312710
rect 575187 312676 575199 312710
rect 575141 312642 575199 312676
rect 575141 312608 575153 312642
rect 575187 312608 575199 312642
rect 575141 312574 575199 312608
rect 575141 312540 575153 312574
rect 575187 312540 575199 312574
rect 575141 312506 575199 312540
rect 575141 312472 575153 312506
rect 575187 312472 575199 312506
rect 575141 312438 575199 312472
rect 575141 312404 575153 312438
rect 575187 312404 575199 312438
rect 575141 312370 575199 312404
rect 575141 312336 575153 312370
rect 575187 312336 575199 312370
rect 575141 312302 575199 312336
rect 575141 312268 575153 312302
rect 575187 312268 575199 312302
rect 575141 312234 575199 312268
rect 575141 312200 575153 312234
rect 575187 312200 575199 312234
rect 575141 312166 575199 312200
rect 575141 312132 575153 312166
rect 575187 312132 575199 312166
rect 575141 312098 575199 312132
rect 575141 312064 575153 312098
rect 575187 312064 575199 312098
rect 575141 312030 575199 312064
rect 575141 311996 575153 312030
rect 575187 311996 575199 312030
rect 575141 311962 575199 311996
rect 575141 311928 575153 311962
rect 575187 311928 575199 311962
rect 575141 311894 575199 311928
rect 575141 311860 575153 311894
rect 575187 311860 575199 311894
rect 575141 311826 575199 311860
rect 575141 311792 575153 311826
rect 575187 311792 575199 311826
rect 575141 311751 575199 311792
rect 575399 312710 575457 312751
rect 575399 312676 575411 312710
rect 575445 312676 575457 312710
rect 575399 312642 575457 312676
rect 575399 312608 575411 312642
rect 575445 312608 575457 312642
rect 575399 312574 575457 312608
rect 575399 312540 575411 312574
rect 575445 312540 575457 312574
rect 575399 312506 575457 312540
rect 575399 312472 575411 312506
rect 575445 312472 575457 312506
rect 575399 312438 575457 312472
rect 575399 312404 575411 312438
rect 575445 312404 575457 312438
rect 575399 312370 575457 312404
rect 575399 312336 575411 312370
rect 575445 312336 575457 312370
rect 575399 312302 575457 312336
rect 575399 312268 575411 312302
rect 575445 312268 575457 312302
rect 575399 312234 575457 312268
rect 575399 312200 575411 312234
rect 575445 312200 575457 312234
rect 575399 312166 575457 312200
rect 575399 312132 575411 312166
rect 575445 312132 575457 312166
rect 575399 312098 575457 312132
rect 575399 312064 575411 312098
rect 575445 312064 575457 312098
rect 575399 312030 575457 312064
rect 575399 311996 575411 312030
rect 575445 311996 575457 312030
rect 575399 311962 575457 311996
rect 575399 311928 575411 311962
rect 575445 311928 575457 311962
rect 575399 311894 575457 311928
rect 575399 311860 575411 311894
rect 575445 311860 575457 311894
rect 575399 311826 575457 311860
rect 575399 311792 575411 311826
rect 575445 311792 575457 311826
rect 575399 311751 575457 311792
rect 575657 312710 575715 312751
rect 575657 312676 575669 312710
rect 575703 312676 575715 312710
rect 575657 312642 575715 312676
rect 575657 312608 575669 312642
rect 575703 312608 575715 312642
rect 575657 312574 575715 312608
rect 575657 312540 575669 312574
rect 575703 312540 575715 312574
rect 575657 312506 575715 312540
rect 575657 312472 575669 312506
rect 575703 312472 575715 312506
rect 575657 312438 575715 312472
rect 575657 312404 575669 312438
rect 575703 312404 575715 312438
rect 575657 312370 575715 312404
rect 575657 312336 575669 312370
rect 575703 312336 575715 312370
rect 575657 312302 575715 312336
rect 575657 312268 575669 312302
rect 575703 312268 575715 312302
rect 575657 312234 575715 312268
rect 575657 312200 575669 312234
rect 575703 312200 575715 312234
rect 575657 312166 575715 312200
rect 575657 312132 575669 312166
rect 575703 312132 575715 312166
rect 575657 312098 575715 312132
rect 575657 312064 575669 312098
rect 575703 312064 575715 312098
rect 575657 312030 575715 312064
rect 575657 311996 575669 312030
rect 575703 311996 575715 312030
rect 575657 311962 575715 311996
rect 575657 311928 575669 311962
rect 575703 311928 575715 311962
rect 575657 311894 575715 311928
rect 575657 311860 575669 311894
rect 575703 311860 575715 311894
rect 575657 311826 575715 311860
rect 575657 311792 575669 311826
rect 575703 311792 575715 311826
rect 575657 311751 575715 311792
rect 575915 312710 575973 312751
rect 575915 312676 575927 312710
rect 575961 312676 575973 312710
rect 575915 312642 575973 312676
rect 575915 312608 575927 312642
rect 575961 312608 575973 312642
rect 575915 312574 575973 312608
rect 575915 312540 575927 312574
rect 575961 312540 575973 312574
rect 575915 312506 575973 312540
rect 575915 312472 575927 312506
rect 575961 312472 575973 312506
rect 575915 312438 575973 312472
rect 575915 312404 575927 312438
rect 575961 312404 575973 312438
rect 575915 312370 575973 312404
rect 575915 312336 575927 312370
rect 575961 312336 575973 312370
rect 575915 312302 575973 312336
rect 575915 312268 575927 312302
rect 575961 312268 575973 312302
rect 575915 312234 575973 312268
rect 575915 312200 575927 312234
rect 575961 312200 575973 312234
rect 575915 312166 575973 312200
rect 575915 312132 575927 312166
rect 575961 312132 575973 312166
rect 575915 312098 575973 312132
rect 575915 312064 575927 312098
rect 575961 312064 575973 312098
rect 575915 312030 575973 312064
rect 575915 311996 575927 312030
rect 575961 311996 575973 312030
rect 575915 311962 575973 311996
rect 575915 311928 575927 311962
rect 575961 311928 575973 311962
rect 575915 311894 575973 311928
rect 575915 311860 575927 311894
rect 575961 311860 575973 311894
rect 575915 311826 575973 311860
rect 575915 311792 575927 311826
rect 575961 311792 575973 311826
rect 575915 311751 575973 311792
rect 576173 312710 576231 312751
rect 576173 312676 576185 312710
rect 576219 312676 576231 312710
rect 576173 312642 576231 312676
rect 576173 312608 576185 312642
rect 576219 312608 576231 312642
rect 576173 312574 576231 312608
rect 576173 312540 576185 312574
rect 576219 312540 576231 312574
rect 576173 312506 576231 312540
rect 576173 312472 576185 312506
rect 576219 312472 576231 312506
rect 576173 312438 576231 312472
rect 576173 312404 576185 312438
rect 576219 312404 576231 312438
rect 576173 312370 576231 312404
rect 576173 312336 576185 312370
rect 576219 312336 576231 312370
rect 576173 312302 576231 312336
rect 576173 312268 576185 312302
rect 576219 312268 576231 312302
rect 576173 312234 576231 312268
rect 576173 312200 576185 312234
rect 576219 312200 576231 312234
rect 576173 312166 576231 312200
rect 576173 312132 576185 312166
rect 576219 312132 576231 312166
rect 576173 312098 576231 312132
rect 576173 312064 576185 312098
rect 576219 312064 576231 312098
rect 576173 312030 576231 312064
rect 576173 311996 576185 312030
rect 576219 311996 576231 312030
rect 576173 311962 576231 311996
rect 576173 311928 576185 311962
rect 576219 311928 576231 311962
rect 576173 311894 576231 311928
rect 576173 311860 576185 311894
rect 576219 311860 576231 311894
rect 576173 311826 576231 311860
rect 576173 311792 576185 311826
rect 576219 311792 576231 311826
rect 576173 311751 576231 311792
rect 576431 312710 576489 312751
rect 576431 312676 576443 312710
rect 576477 312676 576489 312710
rect 576431 312642 576489 312676
rect 576431 312608 576443 312642
rect 576477 312608 576489 312642
rect 576431 312574 576489 312608
rect 576431 312540 576443 312574
rect 576477 312540 576489 312574
rect 576431 312506 576489 312540
rect 576431 312472 576443 312506
rect 576477 312472 576489 312506
rect 576431 312438 576489 312472
rect 576431 312404 576443 312438
rect 576477 312404 576489 312438
rect 576431 312370 576489 312404
rect 576431 312336 576443 312370
rect 576477 312336 576489 312370
rect 576431 312302 576489 312336
rect 576431 312268 576443 312302
rect 576477 312268 576489 312302
rect 576431 312234 576489 312268
rect 576431 312200 576443 312234
rect 576477 312200 576489 312234
rect 576431 312166 576489 312200
rect 576431 312132 576443 312166
rect 576477 312132 576489 312166
rect 576431 312098 576489 312132
rect 576431 312064 576443 312098
rect 576477 312064 576489 312098
rect 576431 312030 576489 312064
rect 576431 311996 576443 312030
rect 576477 311996 576489 312030
rect 576431 311962 576489 311996
rect 576431 311928 576443 311962
rect 576477 311928 576489 311962
rect 576431 311894 576489 311928
rect 576431 311860 576443 311894
rect 576477 311860 576489 311894
rect 576431 311826 576489 311860
rect 576431 311792 576443 311826
rect 576477 311792 576489 311826
rect 576431 311751 576489 311792
rect 576689 312710 576747 312751
rect 576689 312676 576701 312710
rect 576735 312676 576747 312710
rect 576689 312642 576747 312676
rect 576689 312608 576701 312642
rect 576735 312608 576747 312642
rect 576689 312574 576747 312608
rect 576689 312540 576701 312574
rect 576735 312540 576747 312574
rect 576689 312506 576747 312540
rect 576689 312472 576701 312506
rect 576735 312472 576747 312506
rect 576689 312438 576747 312472
rect 576689 312404 576701 312438
rect 576735 312404 576747 312438
rect 576689 312370 576747 312404
rect 576689 312336 576701 312370
rect 576735 312336 576747 312370
rect 576689 312302 576747 312336
rect 576689 312268 576701 312302
rect 576735 312268 576747 312302
rect 576689 312234 576747 312268
rect 576689 312200 576701 312234
rect 576735 312200 576747 312234
rect 576689 312166 576747 312200
rect 576689 312132 576701 312166
rect 576735 312132 576747 312166
rect 576689 312098 576747 312132
rect 576689 312064 576701 312098
rect 576735 312064 576747 312098
rect 576689 312030 576747 312064
rect 576689 311996 576701 312030
rect 576735 311996 576747 312030
rect 576689 311962 576747 311996
rect 576689 311928 576701 311962
rect 576735 311928 576747 311962
rect 576689 311894 576747 311928
rect 576689 311860 576701 311894
rect 576735 311860 576747 311894
rect 576689 311826 576747 311860
rect 576689 311792 576701 311826
rect 576735 311792 576747 311826
rect 576689 311751 576747 311792
rect 576947 312710 577005 312751
rect 576947 312676 576959 312710
rect 576993 312676 577005 312710
rect 576947 312642 577005 312676
rect 576947 312608 576959 312642
rect 576993 312608 577005 312642
rect 576947 312574 577005 312608
rect 576947 312540 576959 312574
rect 576993 312540 577005 312574
rect 576947 312506 577005 312540
rect 576947 312472 576959 312506
rect 576993 312472 577005 312506
rect 576947 312438 577005 312472
rect 576947 312404 576959 312438
rect 576993 312404 577005 312438
rect 576947 312370 577005 312404
rect 576947 312336 576959 312370
rect 576993 312336 577005 312370
rect 576947 312302 577005 312336
rect 576947 312268 576959 312302
rect 576993 312268 577005 312302
rect 576947 312234 577005 312268
rect 576947 312200 576959 312234
rect 576993 312200 577005 312234
rect 576947 312166 577005 312200
rect 576947 312132 576959 312166
rect 576993 312132 577005 312166
rect 576947 312098 577005 312132
rect 576947 312064 576959 312098
rect 576993 312064 577005 312098
rect 576947 312030 577005 312064
rect 576947 311996 576959 312030
rect 576993 311996 577005 312030
rect 576947 311962 577005 311996
rect 576947 311928 576959 311962
rect 576993 311928 577005 311962
rect 576947 311894 577005 311928
rect 576947 311860 576959 311894
rect 576993 311860 577005 311894
rect 576947 311826 577005 311860
rect 576947 311792 576959 311826
rect 576993 311792 577005 311826
rect 576947 311751 577005 311792
rect 577205 312710 577263 312751
rect 577205 312676 577217 312710
rect 577251 312676 577263 312710
rect 577205 312642 577263 312676
rect 577205 312608 577217 312642
rect 577251 312608 577263 312642
rect 577205 312574 577263 312608
rect 577205 312540 577217 312574
rect 577251 312540 577263 312574
rect 577205 312506 577263 312540
rect 577205 312472 577217 312506
rect 577251 312472 577263 312506
rect 577205 312438 577263 312472
rect 577205 312404 577217 312438
rect 577251 312404 577263 312438
rect 577205 312370 577263 312404
rect 577205 312336 577217 312370
rect 577251 312336 577263 312370
rect 577205 312302 577263 312336
rect 577205 312268 577217 312302
rect 577251 312268 577263 312302
rect 577205 312234 577263 312268
rect 577205 312200 577217 312234
rect 577251 312200 577263 312234
rect 577205 312166 577263 312200
rect 577205 312132 577217 312166
rect 577251 312132 577263 312166
rect 577205 312098 577263 312132
rect 577205 312064 577217 312098
rect 577251 312064 577263 312098
rect 577205 312030 577263 312064
rect 577205 311996 577217 312030
rect 577251 311996 577263 312030
rect 577205 311962 577263 311996
rect 577205 311928 577217 311962
rect 577251 311928 577263 311962
rect 577205 311894 577263 311928
rect 577205 311860 577217 311894
rect 577251 311860 577263 311894
rect 577205 311826 577263 311860
rect 577205 311792 577217 311826
rect 577251 311792 577263 311826
rect 577205 311751 577263 311792
rect 577463 312710 577521 312751
rect 577463 312676 577475 312710
rect 577509 312676 577521 312710
rect 577463 312642 577521 312676
rect 577463 312608 577475 312642
rect 577509 312608 577521 312642
rect 577463 312574 577521 312608
rect 577463 312540 577475 312574
rect 577509 312540 577521 312574
rect 577463 312506 577521 312540
rect 577463 312472 577475 312506
rect 577509 312472 577521 312506
rect 577463 312438 577521 312472
rect 577463 312404 577475 312438
rect 577509 312404 577521 312438
rect 577463 312370 577521 312404
rect 577463 312336 577475 312370
rect 577509 312336 577521 312370
rect 577463 312302 577521 312336
rect 577463 312268 577475 312302
rect 577509 312268 577521 312302
rect 577463 312234 577521 312268
rect 577463 312200 577475 312234
rect 577509 312200 577521 312234
rect 577463 312166 577521 312200
rect 577463 312132 577475 312166
rect 577509 312132 577521 312166
rect 577463 312098 577521 312132
rect 577463 312064 577475 312098
rect 577509 312064 577521 312098
rect 577463 312030 577521 312064
rect 577463 311996 577475 312030
rect 577509 311996 577521 312030
rect 577463 311962 577521 311996
rect 577463 311928 577475 311962
rect 577509 311928 577521 311962
rect 577463 311894 577521 311928
rect 577463 311860 577475 311894
rect 577509 311860 577521 311894
rect 577463 311826 577521 311860
rect 577463 311792 577475 311826
rect 577509 311792 577521 311826
rect 577463 311751 577521 311792
rect 577721 312710 577779 312751
rect 577721 312676 577733 312710
rect 577767 312676 577779 312710
rect 577721 312642 577779 312676
rect 577721 312608 577733 312642
rect 577767 312608 577779 312642
rect 577721 312574 577779 312608
rect 577721 312540 577733 312574
rect 577767 312540 577779 312574
rect 577721 312506 577779 312540
rect 577721 312472 577733 312506
rect 577767 312472 577779 312506
rect 577721 312438 577779 312472
rect 577721 312404 577733 312438
rect 577767 312404 577779 312438
rect 577721 312370 577779 312404
rect 577721 312336 577733 312370
rect 577767 312336 577779 312370
rect 577721 312302 577779 312336
rect 577721 312268 577733 312302
rect 577767 312268 577779 312302
rect 577721 312234 577779 312268
rect 577721 312200 577733 312234
rect 577767 312200 577779 312234
rect 577721 312166 577779 312200
rect 577721 312132 577733 312166
rect 577767 312132 577779 312166
rect 577721 312098 577779 312132
rect 577721 312064 577733 312098
rect 577767 312064 577779 312098
rect 577721 312030 577779 312064
rect 577721 311996 577733 312030
rect 577767 311996 577779 312030
rect 577721 311962 577779 311996
rect 577721 311928 577733 311962
rect 577767 311928 577779 311962
rect 577721 311894 577779 311928
rect 577721 311860 577733 311894
rect 577767 311860 577779 311894
rect 577721 311826 577779 311860
rect 577721 311792 577733 311826
rect 577767 311792 577779 311826
rect 577721 311751 577779 311792
rect 577979 312710 578037 312751
rect 577979 312676 577991 312710
rect 578025 312676 578037 312710
rect 577979 312642 578037 312676
rect 577979 312608 577991 312642
rect 578025 312608 578037 312642
rect 577979 312574 578037 312608
rect 577979 312540 577991 312574
rect 578025 312540 578037 312574
rect 577979 312506 578037 312540
rect 577979 312472 577991 312506
rect 578025 312472 578037 312506
rect 577979 312438 578037 312472
rect 577979 312404 577991 312438
rect 578025 312404 578037 312438
rect 577979 312370 578037 312404
rect 577979 312336 577991 312370
rect 578025 312336 578037 312370
rect 577979 312302 578037 312336
rect 577979 312268 577991 312302
rect 578025 312268 578037 312302
rect 577979 312234 578037 312268
rect 577979 312200 577991 312234
rect 578025 312200 578037 312234
rect 577979 312166 578037 312200
rect 577979 312132 577991 312166
rect 578025 312132 578037 312166
rect 577979 312098 578037 312132
rect 577979 312064 577991 312098
rect 578025 312064 578037 312098
rect 577979 312030 578037 312064
rect 577979 311996 577991 312030
rect 578025 311996 578037 312030
rect 577979 311962 578037 311996
rect 577979 311928 577991 311962
rect 578025 311928 578037 311962
rect 577979 311894 578037 311928
rect 577979 311860 577991 311894
rect 578025 311860 578037 311894
rect 577979 311826 578037 311860
rect 577979 311792 577991 311826
rect 578025 311792 578037 311826
rect 577979 311751 578037 311792
rect 578237 312710 578295 312751
rect 578237 312676 578249 312710
rect 578283 312676 578295 312710
rect 578237 312642 578295 312676
rect 578237 312608 578249 312642
rect 578283 312608 578295 312642
rect 578237 312574 578295 312608
rect 578237 312540 578249 312574
rect 578283 312540 578295 312574
rect 578237 312506 578295 312540
rect 578237 312472 578249 312506
rect 578283 312472 578295 312506
rect 578237 312438 578295 312472
rect 578237 312404 578249 312438
rect 578283 312404 578295 312438
rect 578237 312370 578295 312404
rect 578237 312336 578249 312370
rect 578283 312336 578295 312370
rect 578237 312302 578295 312336
rect 578237 312268 578249 312302
rect 578283 312268 578295 312302
rect 578237 312234 578295 312268
rect 578237 312200 578249 312234
rect 578283 312200 578295 312234
rect 578237 312166 578295 312200
rect 578237 312132 578249 312166
rect 578283 312132 578295 312166
rect 578237 312098 578295 312132
rect 578237 312064 578249 312098
rect 578283 312064 578295 312098
rect 578237 312030 578295 312064
rect 578237 311996 578249 312030
rect 578283 311996 578295 312030
rect 578237 311962 578295 311996
rect 578237 311928 578249 311962
rect 578283 311928 578295 311962
rect 578237 311894 578295 311928
rect 578237 311860 578249 311894
rect 578283 311860 578295 311894
rect 578237 311826 578295 311860
rect 578237 311792 578249 311826
rect 578283 311792 578295 311826
rect 578237 311751 578295 311792
rect 578495 312710 578553 312751
rect 578495 312676 578507 312710
rect 578541 312676 578553 312710
rect 578495 312642 578553 312676
rect 578495 312608 578507 312642
rect 578541 312608 578553 312642
rect 578495 312574 578553 312608
rect 578495 312540 578507 312574
rect 578541 312540 578553 312574
rect 578495 312506 578553 312540
rect 578495 312472 578507 312506
rect 578541 312472 578553 312506
rect 578495 312438 578553 312472
rect 578495 312404 578507 312438
rect 578541 312404 578553 312438
rect 578495 312370 578553 312404
rect 578495 312336 578507 312370
rect 578541 312336 578553 312370
rect 578495 312302 578553 312336
rect 578495 312268 578507 312302
rect 578541 312268 578553 312302
rect 578495 312234 578553 312268
rect 578495 312200 578507 312234
rect 578541 312200 578553 312234
rect 578495 312166 578553 312200
rect 578495 312132 578507 312166
rect 578541 312132 578553 312166
rect 578495 312098 578553 312132
rect 578495 312064 578507 312098
rect 578541 312064 578553 312098
rect 578495 312030 578553 312064
rect 578495 311996 578507 312030
rect 578541 311996 578553 312030
rect 578495 311962 578553 311996
rect 578495 311928 578507 311962
rect 578541 311928 578553 311962
rect 578495 311894 578553 311928
rect 578495 311860 578507 311894
rect 578541 311860 578553 311894
rect 578495 311826 578553 311860
rect 578495 311792 578507 311826
rect 578541 311792 578553 311826
rect 578495 311751 578553 311792
rect 578753 312710 578811 312751
rect 578753 312676 578765 312710
rect 578799 312676 578811 312710
rect 578753 312642 578811 312676
rect 578753 312608 578765 312642
rect 578799 312608 578811 312642
rect 578753 312574 578811 312608
rect 578753 312540 578765 312574
rect 578799 312540 578811 312574
rect 578753 312506 578811 312540
rect 578753 312472 578765 312506
rect 578799 312472 578811 312506
rect 578753 312438 578811 312472
rect 578753 312404 578765 312438
rect 578799 312404 578811 312438
rect 578753 312370 578811 312404
rect 578753 312336 578765 312370
rect 578799 312336 578811 312370
rect 578753 312302 578811 312336
rect 578753 312268 578765 312302
rect 578799 312268 578811 312302
rect 578753 312234 578811 312268
rect 578753 312200 578765 312234
rect 578799 312200 578811 312234
rect 578753 312166 578811 312200
rect 578753 312132 578765 312166
rect 578799 312132 578811 312166
rect 578753 312098 578811 312132
rect 578753 312064 578765 312098
rect 578799 312064 578811 312098
rect 578753 312030 578811 312064
rect 578753 311996 578765 312030
rect 578799 311996 578811 312030
rect 578753 311962 578811 311996
rect 578753 311928 578765 311962
rect 578799 311928 578811 311962
rect 578753 311894 578811 311928
rect 578753 311860 578765 311894
rect 578799 311860 578811 311894
rect 578753 311826 578811 311860
rect 578753 311792 578765 311826
rect 578799 311792 578811 311826
rect 578753 311751 578811 311792
rect 579011 312710 579069 312751
rect 579011 312676 579023 312710
rect 579057 312676 579069 312710
rect 579011 312642 579069 312676
rect 579011 312608 579023 312642
rect 579057 312608 579069 312642
rect 579011 312574 579069 312608
rect 579011 312540 579023 312574
rect 579057 312540 579069 312574
rect 579011 312506 579069 312540
rect 579011 312472 579023 312506
rect 579057 312472 579069 312506
rect 579011 312438 579069 312472
rect 579011 312404 579023 312438
rect 579057 312404 579069 312438
rect 579011 312370 579069 312404
rect 579011 312336 579023 312370
rect 579057 312336 579069 312370
rect 579011 312302 579069 312336
rect 579011 312268 579023 312302
rect 579057 312268 579069 312302
rect 579011 312234 579069 312268
rect 579011 312200 579023 312234
rect 579057 312200 579069 312234
rect 579011 312166 579069 312200
rect 579011 312132 579023 312166
rect 579057 312132 579069 312166
rect 579011 312098 579069 312132
rect 579011 312064 579023 312098
rect 579057 312064 579069 312098
rect 579011 312030 579069 312064
rect 579011 311996 579023 312030
rect 579057 311996 579069 312030
rect 579011 311962 579069 311996
rect 579011 311928 579023 311962
rect 579057 311928 579069 311962
rect 579011 311894 579069 311928
rect 579011 311860 579023 311894
rect 579057 311860 579069 311894
rect 579011 311826 579069 311860
rect 579011 311792 579023 311826
rect 579057 311792 579069 311826
rect 579011 311751 579069 311792
rect 579269 312710 579327 312751
rect 579269 312676 579281 312710
rect 579315 312676 579327 312710
rect 579269 312642 579327 312676
rect 579269 312608 579281 312642
rect 579315 312608 579327 312642
rect 579269 312574 579327 312608
rect 579269 312540 579281 312574
rect 579315 312540 579327 312574
rect 579269 312506 579327 312540
rect 579269 312472 579281 312506
rect 579315 312472 579327 312506
rect 579269 312438 579327 312472
rect 579269 312404 579281 312438
rect 579315 312404 579327 312438
rect 579269 312370 579327 312404
rect 579269 312336 579281 312370
rect 579315 312336 579327 312370
rect 579269 312302 579327 312336
rect 579269 312268 579281 312302
rect 579315 312268 579327 312302
rect 579269 312234 579327 312268
rect 579269 312200 579281 312234
rect 579315 312200 579327 312234
rect 579269 312166 579327 312200
rect 579269 312132 579281 312166
rect 579315 312132 579327 312166
rect 579269 312098 579327 312132
rect 579269 312064 579281 312098
rect 579315 312064 579327 312098
rect 579269 312030 579327 312064
rect 579269 311996 579281 312030
rect 579315 311996 579327 312030
rect 579269 311962 579327 311996
rect 579269 311928 579281 311962
rect 579315 311928 579327 311962
rect 579269 311894 579327 311928
rect 579269 311860 579281 311894
rect 579315 311860 579327 311894
rect 579269 311826 579327 311860
rect 579269 311792 579281 311826
rect 579315 311792 579327 311826
rect 579269 311751 579327 311792
rect 579527 312710 579585 312751
rect 579527 312676 579539 312710
rect 579573 312676 579585 312710
rect 579527 312642 579585 312676
rect 579527 312608 579539 312642
rect 579573 312608 579585 312642
rect 579527 312574 579585 312608
rect 579527 312540 579539 312574
rect 579573 312540 579585 312574
rect 579527 312506 579585 312540
rect 579527 312472 579539 312506
rect 579573 312472 579585 312506
rect 579527 312438 579585 312472
rect 579527 312404 579539 312438
rect 579573 312404 579585 312438
rect 579527 312370 579585 312404
rect 579527 312336 579539 312370
rect 579573 312336 579585 312370
rect 579527 312302 579585 312336
rect 579527 312268 579539 312302
rect 579573 312268 579585 312302
rect 579527 312234 579585 312268
rect 579527 312200 579539 312234
rect 579573 312200 579585 312234
rect 579527 312166 579585 312200
rect 579527 312132 579539 312166
rect 579573 312132 579585 312166
rect 579527 312098 579585 312132
rect 579527 312064 579539 312098
rect 579573 312064 579585 312098
rect 579527 312030 579585 312064
rect 579527 311996 579539 312030
rect 579573 311996 579585 312030
rect 579527 311962 579585 311996
rect 579527 311928 579539 311962
rect 579573 311928 579585 311962
rect 579527 311894 579585 311928
rect 579527 311860 579539 311894
rect 579573 311860 579585 311894
rect 579527 311826 579585 311860
rect 579527 311792 579539 311826
rect 579573 311792 579585 311826
rect 579527 311751 579585 311792
rect 579785 312710 579843 312751
rect 579785 312676 579797 312710
rect 579831 312676 579843 312710
rect 579785 312642 579843 312676
rect 579785 312608 579797 312642
rect 579831 312608 579843 312642
rect 579785 312574 579843 312608
rect 579785 312540 579797 312574
rect 579831 312540 579843 312574
rect 579785 312506 579843 312540
rect 579785 312472 579797 312506
rect 579831 312472 579843 312506
rect 579785 312438 579843 312472
rect 579785 312404 579797 312438
rect 579831 312404 579843 312438
rect 579785 312370 579843 312404
rect 579785 312336 579797 312370
rect 579831 312336 579843 312370
rect 579785 312302 579843 312336
rect 579785 312268 579797 312302
rect 579831 312268 579843 312302
rect 579785 312234 579843 312268
rect 579785 312200 579797 312234
rect 579831 312200 579843 312234
rect 579785 312166 579843 312200
rect 579785 312132 579797 312166
rect 579831 312132 579843 312166
rect 579785 312098 579843 312132
rect 579785 312064 579797 312098
rect 579831 312064 579843 312098
rect 579785 312030 579843 312064
rect 579785 311996 579797 312030
rect 579831 311996 579843 312030
rect 579785 311962 579843 311996
rect 579785 311928 579797 311962
rect 579831 311928 579843 311962
rect 579785 311894 579843 311928
rect 579785 311860 579797 311894
rect 579831 311860 579843 311894
rect 579785 311826 579843 311860
rect 579785 311792 579797 311826
rect 579831 311792 579843 311826
rect 579785 311751 579843 311792
rect 580043 312710 580101 312751
rect 580043 312676 580055 312710
rect 580089 312676 580101 312710
rect 580043 312642 580101 312676
rect 580043 312608 580055 312642
rect 580089 312608 580101 312642
rect 580043 312574 580101 312608
rect 580043 312540 580055 312574
rect 580089 312540 580101 312574
rect 580043 312506 580101 312540
rect 580043 312472 580055 312506
rect 580089 312472 580101 312506
rect 580043 312438 580101 312472
rect 580043 312404 580055 312438
rect 580089 312404 580101 312438
rect 580043 312370 580101 312404
rect 580043 312336 580055 312370
rect 580089 312336 580101 312370
rect 580043 312302 580101 312336
rect 580043 312268 580055 312302
rect 580089 312268 580101 312302
rect 580043 312234 580101 312268
rect 580043 312200 580055 312234
rect 580089 312200 580101 312234
rect 580043 312166 580101 312200
rect 580043 312132 580055 312166
rect 580089 312132 580101 312166
rect 580043 312098 580101 312132
rect 580043 312064 580055 312098
rect 580089 312064 580101 312098
rect 580043 312030 580101 312064
rect 580043 311996 580055 312030
rect 580089 311996 580101 312030
rect 580043 311962 580101 311996
rect 580043 311928 580055 311962
rect 580089 311928 580101 311962
rect 580043 311894 580101 311928
rect 580043 311860 580055 311894
rect 580089 311860 580101 311894
rect 580043 311826 580101 311860
rect 580043 311792 580055 311826
rect 580089 311792 580101 311826
rect 580043 311751 580101 311792
rect 580301 312710 580359 312751
rect 580301 312676 580313 312710
rect 580347 312676 580359 312710
rect 580301 312642 580359 312676
rect 580301 312608 580313 312642
rect 580347 312608 580359 312642
rect 580301 312574 580359 312608
rect 580301 312540 580313 312574
rect 580347 312540 580359 312574
rect 580301 312506 580359 312540
rect 580301 312472 580313 312506
rect 580347 312472 580359 312506
rect 580301 312438 580359 312472
rect 580301 312404 580313 312438
rect 580347 312404 580359 312438
rect 580301 312370 580359 312404
rect 580301 312336 580313 312370
rect 580347 312336 580359 312370
rect 580301 312302 580359 312336
rect 580301 312268 580313 312302
rect 580347 312268 580359 312302
rect 580301 312234 580359 312268
rect 580301 312200 580313 312234
rect 580347 312200 580359 312234
rect 580301 312166 580359 312200
rect 580301 312132 580313 312166
rect 580347 312132 580359 312166
rect 580301 312098 580359 312132
rect 580301 312064 580313 312098
rect 580347 312064 580359 312098
rect 580301 312030 580359 312064
rect 580301 311996 580313 312030
rect 580347 311996 580359 312030
rect 580301 311962 580359 311996
rect 580301 311928 580313 311962
rect 580347 311928 580359 311962
rect 580301 311894 580359 311928
rect 580301 311860 580313 311894
rect 580347 311860 580359 311894
rect 580301 311826 580359 311860
rect 580301 311792 580313 311826
rect 580347 311792 580359 311826
rect 580301 311751 580359 311792
<< ndiffc >>
rect 560675 493374 560709 493408
rect 560675 493306 560709 493340
rect 560675 493238 560709 493272
rect 560675 493170 560709 493204
rect 560675 493102 560709 493136
rect 560675 493034 560709 493068
rect 560675 492966 560709 493000
rect 560675 492898 560709 492932
rect 560675 492830 560709 492864
rect 560675 492762 560709 492796
rect 560675 492694 560709 492728
rect 560675 492626 560709 492660
rect 560675 492558 560709 492592
rect 560675 492490 560709 492524
rect 560933 493374 560967 493408
rect 560933 493306 560967 493340
rect 560933 493238 560967 493272
rect 560933 493170 560967 493204
rect 560933 493102 560967 493136
rect 560933 493034 560967 493068
rect 560933 492966 560967 493000
rect 560933 492898 560967 492932
rect 560933 492830 560967 492864
rect 560933 492762 560967 492796
rect 560933 492694 560967 492728
rect 560933 492626 560967 492660
rect 560933 492558 560967 492592
rect 560933 492490 560967 492524
rect 561191 493374 561225 493408
rect 561191 493306 561225 493340
rect 561191 493238 561225 493272
rect 561191 493170 561225 493204
rect 561191 493102 561225 493136
rect 561191 493034 561225 493068
rect 561191 492966 561225 493000
rect 561191 492898 561225 492932
rect 561191 492830 561225 492864
rect 561191 492762 561225 492796
rect 561191 492694 561225 492728
rect 561191 492626 561225 492660
rect 561191 492558 561225 492592
rect 561191 492490 561225 492524
rect 561449 493374 561483 493408
rect 561449 493306 561483 493340
rect 561449 493238 561483 493272
rect 561449 493170 561483 493204
rect 561449 493102 561483 493136
rect 561449 493034 561483 493068
rect 561449 492966 561483 493000
rect 561449 492898 561483 492932
rect 561449 492830 561483 492864
rect 561449 492762 561483 492796
rect 561449 492694 561483 492728
rect 561449 492626 561483 492660
rect 561449 492558 561483 492592
rect 561449 492490 561483 492524
rect 561707 493374 561741 493408
rect 561707 493306 561741 493340
rect 561707 493238 561741 493272
rect 561707 493170 561741 493204
rect 561707 493102 561741 493136
rect 561707 493034 561741 493068
rect 561707 492966 561741 493000
rect 561707 492898 561741 492932
rect 561707 492830 561741 492864
rect 561707 492762 561741 492796
rect 561707 492694 561741 492728
rect 561707 492626 561741 492660
rect 561707 492558 561741 492592
rect 561707 492490 561741 492524
rect 561965 493374 561999 493408
rect 561965 493306 561999 493340
rect 561965 493238 561999 493272
rect 561965 493170 561999 493204
rect 561965 493102 561999 493136
rect 561965 493034 561999 493068
rect 561965 492966 561999 493000
rect 561965 492898 561999 492932
rect 561965 492830 561999 492864
rect 561965 492762 561999 492796
rect 561965 492694 561999 492728
rect 561965 492626 561999 492660
rect 561965 492558 561999 492592
rect 561965 492490 561999 492524
rect 562223 493374 562257 493408
rect 562223 493306 562257 493340
rect 562223 493238 562257 493272
rect 562223 493170 562257 493204
rect 562223 493102 562257 493136
rect 562223 493034 562257 493068
rect 562223 492966 562257 493000
rect 562223 492898 562257 492932
rect 562223 492830 562257 492864
rect 562223 492762 562257 492796
rect 562223 492694 562257 492728
rect 562223 492626 562257 492660
rect 562223 492558 562257 492592
rect 562223 492490 562257 492524
rect 562481 493374 562515 493408
rect 562481 493306 562515 493340
rect 562481 493238 562515 493272
rect 562481 493170 562515 493204
rect 562481 493102 562515 493136
rect 562481 493034 562515 493068
rect 562481 492966 562515 493000
rect 562481 492898 562515 492932
rect 562481 492830 562515 492864
rect 562481 492762 562515 492796
rect 562481 492694 562515 492728
rect 562481 492626 562515 492660
rect 562481 492558 562515 492592
rect 562481 492490 562515 492524
rect 562739 493374 562773 493408
rect 562739 493306 562773 493340
rect 562739 493238 562773 493272
rect 562739 493170 562773 493204
rect 562739 493102 562773 493136
rect 562739 493034 562773 493068
rect 562739 492966 562773 493000
rect 562739 492898 562773 492932
rect 562739 492830 562773 492864
rect 562739 492762 562773 492796
rect 562739 492694 562773 492728
rect 562739 492626 562773 492660
rect 562739 492558 562773 492592
rect 562739 492490 562773 492524
rect 562997 493374 563031 493408
rect 562997 493306 563031 493340
rect 562997 493238 563031 493272
rect 562997 493170 563031 493204
rect 562997 493102 563031 493136
rect 562997 493034 563031 493068
rect 562997 492966 563031 493000
rect 562997 492898 563031 492932
rect 562997 492830 563031 492864
rect 562997 492762 563031 492796
rect 562997 492694 563031 492728
rect 562997 492626 563031 492660
rect 562997 492558 563031 492592
rect 562997 492490 563031 492524
rect 563255 493374 563289 493408
rect 563255 493306 563289 493340
rect 563255 493238 563289 493272
rect 563255 493170 563289 493204
rect 563255 493102 563289 493136
rect 563255 493034 563289 493068
rect 563255 492966 563289 493000
rect 563255 492898 563289 492932
rect 563255 492830 563289 492864
rect 563255 492762 563289 492796
rect 563255 492694 563289 492728
rect 563255 492626 563289 492660
rect 563255 492558 563289 492592
rect 563255 492490 563289 492524
rect 563513 493374 563547 493408
rect 563513 493306 563547 493340
rect 563513 493238 563547 493272
rect 563513 493170 563547 493204
rect 563513 493102 563547 493136
rect 563513 493034 563547 493068
rect 563513 492966 563547 493000
rect 563513 492898 563547 492932
rect 563513 492830 563547 492864
rect 563513 492762 563547 492796
rect 563513 492694 563547 492728
rect 563513 492626 563547 492660
rect 563513 492558 563547 492592
rect 563513 492490 563547 492524
rect 563771 493374 563805 493408
rect 563771 493306 563805 493340
rect 563771 493238 563805 493272
rect 563771 493170 563805 493204
rect 563771 493102 563805 493136
rect 563771 493034 563805 493068
rect 563771 492966 563805 493000
rect 563771 492898 563805 492932
rect 563771 492830 563805 492864
rect 563771 492762 563805 492796
rect 563771 492694 563805 492728
rect 563771 492626 563805 492660
rect 563771 492558 563805 492592
rect 563771 492490 563805 492524
rect 564029 493374 564063 493408
rect 564029 493306 564063 493340
rect 564029 493238 564063 493272
rect 564029 493170 564063 493204
rect 564029 493102 564063 493136
rect 564029 493034 564063 493068
rect 564029 492966 564063 493000
rect 564029 492898 564063 492932
rect 564029 492830 564063 492864
rect 564029 492762 564063 492796
rect 564029 492694 564063 492728
rect 564029 492626 564063 492660
rect 564029 492558 564063 492592
rect 564029 492490 564063 492524
rect 564287 493374 564321 493408
rect 564287 493306 564321 493340
rect 564287 493238 564321 493272
rect 564287 493170 564321 493204
rect 564287 493102 564321 493136
rect 564287 493034 564321 493068
rect 564287 492966 564321 493000
rect 564287 492898 564321 492932
rect 564287 492830 564321 492864
rect 564287 492762 564321 492796
rect 564287 492694 564321 492728
rect 564287 492626 564321 492660
rect 564287 492558 564321 492592
rect 564287 492490 564321 492524
rect 564545 493374 564579 493408
rect 564545 493306 564579 493340
rect 564545 493238 564579 493272
rect 564545 493170 564579 493204
rect 564545 493102 564579 493136
rect 564545 493034 564579 493068
rect 564545 492966 564579 493000
rect 564545 492898 564579 492932
rect 564545 492830 564579 492864
rect 564545 492762 564579 492796
rect 564545 492694 564579 492728
rect 564545 492626 564579 492660
rect 564545 492558 564579 492592
rect 564545 492490 564579 492524
rect 564803 493374 564837 493408
rect 564803 493306 564837 493340
rect 564803 493238 564837 493272
rect 564803 493170 564837 493204
rect 564803 493102 564837 493136
rect 564803 493034 564837 493068
rect 564803 492966 564837 493000
rect 564803 492898 564837 492932
rect 564803 492830 564837 492864
rect 564803 492762 564837 492796
rect 564803 492694 564837 492728
rect 564803 492626 564837 492660
rect 564803 492558 564837 492592
rect 564803 492490 564837 492524
rect 565061 493374 565095 493408
rect 565061 493306 565095 493340
rect 565061 493238 565095 493272
rect 565061 493170 565095 493204
rect 565061 493102 565095 493136
rect 565061 493034 565095 493068
rect 565061 492966 565095 493000
rect 565061 492898 565095 492932
rect 565061 492830 565095 492864
rect 565061 492762 565095 492796
rect 565061 492694 565095 492728
rect 565061 492626 565095 492660
rect 565061 492558 565095 492592
rect 565061 492490 565095 492524
rect 565319 493374 565353 493408
rect 565319 493306 565353 493340
rect 565319 493238 565353 493272
rect 565319 493170 565353 493204
rect 565319 493102 565353 493136
rect 565319 493034 565353 493068
rect 565319 492966 565353 493000
rect 565319 492898 565353 492932
rect 565319 492830 565353 492864
rect 565319 492762 565353 492796
rect 565319 492694 565353 492728
rect 565319 492626 565353 492660
rect 565319 492558 565353 492592
rect 565319 492490 565353 492524
rect 565577 493374 565611 493408
rect 565577 493306 565611 493340
rect 565577 493238 565611 493272
rect 565577 493170 565611 493204
rect 565577 493102 565611 493136
rect 565577 493034 565611 493068
rect 565577 492966 565611 493000
rect 565577 492898 565611 492932
rect 565577 492830 565611 492864
rect 565577 492762 565611 492796
rect 565577 492694 565611 492728
rect 565577 492626 565611 492660
rect 565577 492558 565611 492592
rect 565577 492490 565611 492524
rect 565835 493374 565869 493408
rect 565835 493306 565869 493340
rect 565835 493238 565869 493272
rect 565835 493170 565869 493204
rect 565835 493102 565869 493136
rect 565835 493034 565869 493068
rect 565835 492966 565869 493000
rect 565835 492898 565869 492932
rect 565835 492830 565869 492864
rect 565835 492762 565869 492796
rect 565835 492694 565869 492728
rect 565835 492626 565869 492660
rect 565835 492558 565869 492592
rect 565835 492490 565869 492524
rect 560611 404232 560645 404266
rect 560611 404164 560645 404198
rect 560611 404096 560645 404130
rect 560611 404028 560645 404062
rect 560611 403960 560645 403994
rect 560611 403892 560645 403926
rect 560611 403824 560645 403858
rect 560611 403756 560645 403790
rect 560611 403688 560645 403722
rect 560611 403620 560645 403654
rect 560611 403552 560645 403586
rect 560611 403484 560645 403518
rect 560611 403416 560645 403450
rect 560611 403348 560645 403382
rect 560869 404232 560903 404266
rect 560869 404164 560903 404198
rect 560869 404096 560903 404130
rect 560869 404028 560903 404062
rect 560869 403960 560903 403994
rect 560869 403892 560903 403926
rect 560869 403824 560903 403858
rect 560869 403756 560903 403790
rect 560869 403688 560903 403722
rect 560869 403620 560903 403654
rect 560869 403552 560903 403586
rect 560869 403484 560903 403518
rect 560869 403416 560903 403450
rect 560869 403348 560903 403382
rect 561127 404232 561161 404266
rect 561127 404164 561161 404198
rect 561127 404096 561161 404130
rect 561127 404028 561161 404062
rect 561127 403960 561161 403994
rect 561127 403892 561161 403926
rect 561127 403824 561161 403858
rect 561127 403756 561161 403790
rect 561127 403688 561161 403722
rect 561127 403620 561161 403654
rect 561127 403552 561161 403586
rect 561127 403484 561161 403518
rect 561127 403416 561161 403450
rect 561127 403348 561161 403382
rect 561385 404232 561419 404266
rect 561385 404164 561419 404198
rect 561385 404096 561419 404130
rect 561385 404028 561419 404062
rect 561385 403960 561419 403994
rect 561385 403892 561419 403926
rect 561385 403824 561419 403858
rect 561385 403756 561419 403790
rect 561385 403688 561419 403722
rect 561385 403620 561419 403654
rect 561385 403552 561419 403586
rect 561385 403484 561419 403518
rect 561385 403416 561419 403450
rect 561385 403348 561419 403382
rect 561643 404232 561677 404266
rect 561643 404164 561677 404198
rect 561643 404096 561677 404130
rect 561643 404028 561677 404062
rect 561643 403960 561677 403994
rect 561643 403892 561677 403926
rect 561643 403824 561677 403858
rect 561643 403756 561677 403790
rect 561643 403688 561677 403722
rect 561643 403620 561677 403654
rect 561643 403552 561677 403586
rect 561643 403484 561677 403518
rect 561643 403416 561677 403450
rect 561643 403348 561677 403382
rect 561901 404232 561935 404266
rect 561901 404164 561935 404198
rect 561901 404096 561935 404130
rect 561901 404028 561935 404062
rect 561901 403960 561935 403994
rect 561901 403892 561935 403926
rect 561901 403824 561935 403858
rect 561901 403756 561935 403790
rect 561901 403688 561935 403722
rect 561901 403620 561935 403654
rect 561901 403552 561935 403586
rect 561901 403484 561935 403518
rect 561901 403416 561935 403450
rect 561901 403348 561935 403382
rect 562159 404232 562193 404266
rect 562159 404164 562193 404198
rect 562159 404096 562193 404130
rect 562159 404028 562193 404062
rect 562159 403960 562193 403994
rect 562159 403892 562193 403926
rect 562159 403824 562193 403858
rect 562159 403756 562193 403790
rect 562159 403688 562193 403722
rect 562159 403620 562193 403654
rect 562159 403552 562193 403586
rect 562159 403484 562193 403518
rect 562159 403416 562193 403450
rect 562159 403348 562193 403382
rect 562417 404232 562451 404266
rect 562417 404164 562451 404198
rect 562417 404096 562451 404130
rect 562417 404028 562451 404062
rect 562417 403960 562451 403994
rect 562417 403892 562451 403926
rect 562417 403824 562451 403858
rect 562417 403756 562451 403790
rect 562417 403688 562451 403722
rect 562417 403620 562451 403654
rect 562417 403552 562451 403586
rect 562417 403484 562451 403518
rect 562417 403416 562451 403450
rect 562417 403348 562451 403382
rect 562675 404232 562709 404266
rect 562675 404164 562709 404198
rect 562675 404096 562709 404130
rect 562675 404028 562709 404062
rect 562675 403960 562709 403994
rect 562675 403892 562709 403926
rect 562675 403824 562709 403858
rect 562675 403756 562709 403790
rect 562675 403688 562709 403722
rect 562675 403620 562709 403654
rect 562675 403552 562709 403586
rect 562675 403484 562709 403518
rect 562675 403416 562709 403450
rect 562675 403348 562709 403382
rect 562933 404232 562967 404266
rect 562933 404164 562967 404198
rect 562933 404096 562967 404130
rect 562933 404028 562967 404062
rect 562933 403960 562967 403994
rect 562933 403892 562967 403926
rect 562933 403824 562967 403858
rect 562933 403756 562967 403790
rect 562933 403688 562967 403722
rect 562933 403620 562967 403654
rect 562933 403552 562967 403586
rect 562933 403484 562967 403518
rect 562933 403416 562967 403450
rect 562933 403348 562967 403382
rect 563191 404232 563225 404266
rect 563191 404164 563225 404198
rect 563191 404096 563225 404130
rect 563191 404028 563225 404062
rect 563191 403960 563225 403994
rect 563191 403892 563225 403926
rect 563191 403824 563225 403858
rect 563191 403756 563225 403790
rect 563191 403688 563225 403722
rect 563191 403620 563225 403654
rect 563191 403552 563225 403586
rect 563191 403484 563225 403518
rect 563191 403416 563225 403450
rect 563191 403348 563225 403382
rect 563449 404232 563483 404266
rect 563449 404164 563483 404198
rect 563449 404096 563483 404130
rect 563449 404028 563483 404062
rect 563449 403960 563483 403994
rect 563449 403892 563483 403926
rect 563449 403824 563483 403858
rect 563449 403756 563483 403790
rect 563449 403688 563483 403722
rect 563449 403620 563483 403654
rect 563449 403552 563483 403586
rect 563449 403484 563483 403518
rect 563449 403416 563483 403450
rect 563449 403348 563483 403382
rect 563707 404232 563741 404266
rect 563707 404164 563741 404198
rect 563707 404096 563741 404130
rect 563707 404028 563741 404062
rect 563707 403960 563741 403994
rect 563707 403892 563741 403926
rect 563707 403824 563741 403858
rect 563707 403756 563741 403790
rect 563707 403688 563741 403722
rect 563707 403620 563741 403654
rect 563707 403552 563741 403586
rect 563707 403484 563741 403518
rect 563707 403416 563741 403450
rect 563707 403348 563741 403382
rect 563965 404232 563999 404266
rect 563965 404164 563999 404198
rect 563965 404096 563999 404130
rect 563965 404028 563999 404062
rect 563965 403960 563999 403994
rect 563965 403892 563999 403926
rect 563965 403824 563999 403858
rect 563965 403756 563999 403790
rect 563965 403688 563999 403722
rect 563965 403620 563999 403654
rect 563965 403552 563999 403586
rect 563965 403484 563999 403518
rect 563965 403416 563999 403450
rect 563965 403348 563999 403382
rect 564223 404232 564257 404266
rect 564223 404164 564257 404198
rect 564223 404096 564257 404130
rect 564223 404028 564257 404062
rect 564223 403960 564257 403994
rect 564223 403892 564257 403926
rect 564223 403824 564257 403858
rect 564223 403756 564257 403790
rect 564223 403688 564257 403722
rect 564223 403620 564257 403654
rect 564223 403552 564257 403586
rect 564223 403484 564257 403518
rect 564223 403416 564257 403450
rect 564223 403348 564257 403382
rect 564481 404232 564515 404266
rect 564481 404164 564515 404198
rect 564481 404096 564515 404130
rect 564481 404028 564515 404062
rect 564481 403960 564515 403994
rect 564481 403892 564515 403926
rect 564481 403824 564515 403858
rect 564481 403756 564515 403790
rect 564481 403688 564515 403722
rect 564481 403620 564515 403654
rect 564481 403552 564515 403586
rect 564481 403484 564515 403518
rect 564481 403416 564515 403450
rect 564481 403348 564515 403382
rect 564739 404232 564773 404266
rect 564739 404164 564773 404198
rect 564739 404096 564773 404130
rect 564739 404028 564773 404062
rect 564739 403960 564773 403994
rect 564739 403892 564773 403926
rect 564739 403824 564773 403858
rect 564739 403756 564773 403790
rect 564739 403688 564773 403722
rect 564739 403620 564773 403654
rect 564739 403552 564773 403586
rect 564739 403484 564773 403518
rect 564739 403416 564773 403450
rect 564739 403348 564773 403382
rect 564997 404232 565031 404266
rect 564997 404164 565031 404198
rect 564997 404096 565031 404130
rect 564997 404028 565031 404062
rect 564997 403960 565031 403994
rect 564997 403892 565031 403926
rect 564997 403824 565031 403858
rect 564997 403756 565031 403790
rect 564997 403688 565031 403722
rect 564997 403620 565031 403654
rect 564997 403552 565031 403586
rect 564997 403484 565031 403518
rect 564997 403416 565031 403450
rect 564997 403348 565031 403382
rect 565255 404232 565289 404266
rect 565255 404164 565289 404198
rect 565255 404096 565289 404130
rect 565255 404028 565289 404062
rect 565255 403960 565289 403994
rect 565255 403892 565289 403926
rect 565255 403824 565289 403858
rect 565255 403756 565289 403790
rect 565255 403688 565289 403722
rect 565255 403620 565289 403654
rect 565255 403552 565289 403586
rect 565255 403484 565289 403518
rect 565255 403416 565289 403450
rect 565255 403348 565289 403382
rect 565513 404232 565547 404266
rect 565513 404164 565547 404198
rect 565513 404096 565547 404130
rect 565513 404028 565547 404062
rect 565513 403960 565547 403994
rect 565513 403892 565547 403926
rect 565513 403824 565547 403858
rect 565513 403756 565547 403790
rect 565513 403688 565547 403722
rect 565513 403620 565547 403654
rect 565513 403552 565547 403586
rect 565513 403484 565547 403518
rect 565513 403416 565547 403450
rect 565513 403348 565547 403382
rect 565771 404232 565805 404266
rect 565771 404164 565805 404198
rect 565771 404096 565805 404130
rect 565771 404028 565805 404062
rect 565771 403960 565805 403994
rect 565771 403892 565805 403926
rect 565771 403824 565805 403858
rect 565771 403756 565805 403790
rect 565771 403688 565805 403722
rect 565771 403620 565805 403654
rect 565771 403552 565805 403586
rect 565771 403484 565805 403518
rect 565771 403416 565805 403450
rect 565771 403348 565805 403382
rect 560567 358914 560601 358948
rect 560567 358846 560601 358880
rect 560567 358778 560601 358812
rect 560567 358710 560601 358744
rect 560567 358642 560601 358676
rect 560567 358574 560601 358608
rect 560567 358506 560601 358540
rect 560567 358438 560601 358472
rect 560567 358370 560601 358404
rect 560567 358302 560601 358336
rect 560567 358234 560601 358268
rect 560567 358166 560601 358200
rect 560567 358098 560601 358132
rect 560567 358030 560601 358064
rect 560825 358914 560859 358948
rect 560825 358846 560859 358880
rect 560825 358778 560859 358812
rect 560825 358710 560859 358744
rect 560825 358642 560859 358676
rect 560825 358574 560859 358608
rect 560825 358506 560859 358540
rect 560825 358438 560859 358472
rect 560825 358370 560859 358404
rect 560825 358302 560859 358336
rect 560825 358234 560859 358268
rect 560825 358166 560859 358200
rect 560825 358098 560859 358132
rect 560825 358030 560859 358064
rect 561083 358914 561117 358948
rect 561083 358846 561117 358880
rect 561083 358778 561117 358812
rect 561083 358710 561117 358744
rect 561083 358642 561117 358676
rect 561083 358574 561117 358608
rect 561083 358506 561117 358540
rect 561083 358438 561117 358472
rect 561083 358370 561117 358404
rect 561083 358302 561117 358336
rect 561083 358234 561117 358268
rect 561083 358166 561117 358200
rect 561083 358098 561117 358132
rect 561083 358030 561117 358064
rect 561341 358914 561375 358948
rect 561341 358846 561375 358880
rect 561341 358778 561375 358812
rect 561341 358710 561375 358744
rect 561341 358642 561375 358676
rect 561341 358574 561375 358608
rect 561341 358506 561375 358540
rect 561341 358438 561375 358472
rect 561341 358370 561375 358404
rect 561341 358302 561375 358336
rect 561341 358234 561375 358268
rect 561341 358166 561375 358200
rect 561341 358098 561375 358132
rect 561341 358030 561375 358064
rect 561599 358914 561633 358948
rect 561599 358846 561633 358880
rect 561599 358778 561633 358812
rect 561599 358710 561633 358744
rect 561599 358642 561633 358676
rect 561599 358574 561633 358608
rect 561599 358506 561633 358540
rect 561599 358438 561633 358472
rect 561599 358370 561633 358404
rect 561599 358302 561633 358336
rect 561599 358234 561633 358268
rect 561599 358166 561633 358200
rect 561599 358098 561633 358132
rect 561599 358030 561633 358064
rect 561857 358914 561891 358948
rect 561857 358846 561891 358880
rect 561857 358778 561891 358812
rect 561857 358710 561891 358744
rect 561857 358642 561891 358676
rect 561857 358574 561891 358608
rect 561857 358506 561891 358540
rect 561857 358438 561891 358472
rect 561857 358370 561891 358404
rect 561857 358302 561891 358336
rect 561857 358234 561891 358268
rect 561857 358166 561891 358200
rect 561857 358098 561891 358132
rect 561857 358030 561891 358064
rect 562115 358914 562149 358948
rect 562115 358846 562149 358880
rect 562115 358778 562149 358812
rect 562115 358710 562149 358744
rect 562115 358642 562149 358676
rect 562115 358574 562149 358608
rect 562115 358506 562149 358540
rect 562115 358438 562149 358472
rect 562115 358370 562149 358404
rect 562115 358302 562149 358336
rect 562115 358234 562149 358268
rect 562115 358166 562149 358200
rect 562115 358098 562149 358132
rect 562115 358030 562149 358064
rect 562373 358914 562407 358948
rect 562373 358846 562407 358880
rect 562373 358778 562407 358812
rect 562373 358710 562407 358744
rect 562373 358642 562407 358676
rect 562373 358574 562407 358608
rect 562373 358506 562407 358540
rect 562373 358438 562407 358472
rect 562373 358370 562407 358404
rect 562373 358302 562407 358336
rect 562373 358234 562407 358268
rect 562373 358166 562407 358200
rect 562373 358098 562407 358132
rect 562373 358030 562407 358064
rect 562631 358914 562665 358948
rect 562631 358846 562665 358880
rect 562631 358778 562665 358812
rect 562631 358710 562665 358744
rect 562631 358642 562665 358676
rect 562631 358574 562665 358608
rect 562631 358506 562665 358540
rect 562631 358438 562665 358472
rect 562631 358370 562665 358404
rect 562631 358302 562665 358336
rect 562631 358234 562665 358268
rect 562631 358166 562665 358200
rect 562631 358098 562665 358132
rect 562631 358030 562665 358064
rect 562889 358914 562923 358948
rect 562889 358846 562923 358880
rect 562889 358778 562923 358812
rect 562889 358710 562923 358744
rect 562889 358642 562923 358676
rect 562889 358574 562923 358608
rect 562889 358506 562923 358540
rect 562889 358438 562923 358472
rect 562889 358370 562923 358404
rect 562889 358302 562923 358336
rect 562889 358234 562923 358268
rect 562889 358166 562923 358200
rect 562889 358098 562923 358132
rect 562889 358030 562923 358064
rect 563147 358914 563181 358948
rect 563147 358846 563181 358880
rect 563147 358778 563181 358812
rect 563147 358710 563181 358744
rect 563147 358642 563181 358676
rect 563147 358574 563181 358608
rect 563147 358506 563181 358540
rect 563147 358438 563181 358472
rect 563147 358370 563181 358404
rect 563147 358302 563181 358336
rect 563147 358234 563181 358268
rect 563147 358166 563181 358200
rect 563147 358098 563181 358132
rect 563147 358030 563181 358064
rect 563405 358914 563439 358948
rect 563405 358846 563439 358880
rect 563405 358778 563439 358812
rect 563405 358710 563439 358744
rect 563405 358642 563439 358676
rect 563405 358574 563439 358608
rect 563405 358506 563439 358540
rect 563405 358438 563439 358472
rect 563405 358370 563439 358404
rect 563405 358302 563439 358336
rect 563405 358234 563439 358268
rect 563405 358166 563439 358200
rect 563405 358098 563439 358132
rect 563405 358030 563439 358064
rect 563663 358914 563697 358948
rect 563663 358846 563697 358880
rect 563663 358778 563697 358812
rect 563663 358710 563697 358744
rect 563663 358642 563697 358676
rect 563663 358574 563697 358608
rect 563663 358506 563697 358540
rect 563663 358438 563697 358472
rect 563663 358370 563697 358404
rect 563663 358302 563697 358336
rect 563663 358234 563697 358268
rect 563663 358166 563697 358200
rect 563663 358098 563697 358132
rect 563663 358030 563697 358064
rect 563921 358914 563955 358948
rect 563921 358846 563955 358880
rect 563921 358778 563955 358812
rect 563921 358710 563955 358744
rect 563921 358642 563955 358676
rect 563921 358574 563955 358608
rect 563921 358506 563955 358540
rect 563921 358438 563955 358472
rect 563921 358370 563955 358404
rect 563921 358302 563955 358336
rect 563921 358234 563955 358268
rect 563921 358166 563955 358200
rect 563921 358098 563955 358132
rect 563921 358030 563955 358064
rect 564179 358914 564213 358948
rect 564179 358846 564213 358880
rect 564179 358778 564213 358812
rect 564179 358710 564213 358744
rect 564179 358642 564213 358676
rect 564179 358574 564213 358608
rect 564179 358506 564213 358540
rect 564179 358438 564213 358472
rect 564179 358370 564213 358404
rect 564179 358302 564213 358336
rect 564179 358234 564213 358268
rect 564179 358166 564213 358200
rect 564179 358098 564213 358132
rect 564179 358030 564213 358064
rect 564437 358914 564471 358948
rect 564437 358846 564471 358880
rect 564437 358778 564471 358812
rect 564437 358710 564471 358744
rect 564437 358642 564471 358676
rect 564437 358574 564471 358608
rect 564437 358506 564471 358540
rect 564437 358438 564471 358472
rect 564437 358370 564471 358404
rect 564437 358302 564471 358336
rect 564437 358234 564471 358268
rect 564437 358166 564471 358200
rect 564437 358098 564471 358132
rect 564437 358030 564471 358064
rect 564695 358914 564729 358948
rect 564695 358846 564729 358880
rect 564695 358778 564729 358812
rect 564695 358710 564729 358744
rect 564695 358642 564729 358676
rect 564695 358574 564729 358608
rect 564695 358506 564729 358540
rect 564695 358438 564729 358472
rect 564695 358370 564729 358404
rect 564695 358302 564729 358336
rect 564695 358234 564729 358268
rect 564695 358166 564729 358200
rect 564695 358098 564729 358132
rect 564695 358030 564729 358064
rect 564953 358914 564987 358948
rect 564953 358846 564987 358880
rect 564953 358778 564987 358812
rect 564953 358710 564987 358744
rect 564953 358642 564987 358676
rect 564953 358574 564987 358608
rect 564953 358506 564987 358540
rect 564953 358438 564987 358472
rect 564953 358370 564987 358404
rect 564953 358302 564987 358336
rect 564953 358234 564987 358268
rect 564953 358166 564987 358200
rect 564953 358098 564987 358132
rect 564953 358030 564987 358064
rect 565211 358914 565245 358948
rect 565211 358846 565245 358880
rect 565211 358778 565245 358812
rect 565211 358710 565245 358744
rect 565211 358642 565245 358676
rect 565211 358574 565245 358608
rect 565211 358506 565245 358540
rect 565211 358438 565245 358472
rect 565211 358370 565245 358404
rect 565211 358302 565245 358336
rect 565211 358234 565245 358268
rect 565211 358166 565245 358200
rect 565211 358098 565245 358132
rect 565211 358030 565245 358064
rect 565469 358914 565503 358948
rect 565469 358846 565503 358880
rect 565469 358778 565503 358812
rect 565469 358710 565503 358744
rect 565469 358642 565503 358676
rect 565469 358574 565503 358608
rect 565469 358506 565503 358540
rect 565469 358438 565503 358472
rect 565469 358370 565503 358404
rect 565469 358302 565503 358336
rect 565469 358234 565503 358268
rect 565469 358166 565503 358200
rect 565469 358098 565503 358132
rect 565469 358030 565503 358064
rect 565727 358914 565761 358948
rect 565727 358846 565761 358880
rect 565727 358778 565761 358812
rect 565727 358710 565761 358744
rect 565727 358642 565761 358676
rect 565727 358574 565761 358608
rect 565727 358506 565761 358540
rect 565727 358438 565761 358472
rect 565727 358370 565761 358404
rect 565727 358302 565761 358336
rect 565727 358234 565761 358268
rect 565727 358166 565761 358200
rect 565727 358098 565761 358132
rect 565727 358030 565761 358064
rect 560429 312606 560463 312640
rect 560429 312538 560463 312572
rect 560429 312470 560463 312504
rect 560429 312402 560463 312436
rect 560429 312334 560463 312368
rect 560429 312266 560463 312300
rect 560429 312198 560463 312232
rect 560429 312130 560463 312164
rect 560429 312062 560463 312096
rect 560429 311994 560463 312028
rect 560429 311926 560463 311960
rect 560429 311858 560463 311892
rect 560429 311790 560463 311824
rect 560429 311722 560463 311756
rect 560687 312606 560721 312640
rect 560687 312538 560721 312572
rect 560687 312470 560721 312504
rect 560687 312402 560721 312436
rect 560687 312334 560721 312368
rect 560687 312266 560721 312300
rect 560687 312198 560721 312232
rect 560687 312130 560721 312164
rect 560687 312062 560721 312096
rect 560687 311994 560721 312028
rect 560687 311926 560721 311960
rect 560687 311858 560721 311892
rect 560687 311790 560721 311824
rect 560687 311722 560721 311756
rect 560945 312606 560979 312640
rect 560945 312538 560979 312572
rect 560945 312470 560979 312504
rect 560945 312402 560979 312436
rect 560945 312334 560979 312368
rect 560945 312266 560979 312300
rect 560945 312198 560979 312232
rect 560945 312130 560979 312164
rect 560945 312062 560979 312096
rect 560945 311994 560979 312028
rect 560945 311926 560979 311960
rect 560945 311858 560979 311892
rect 560945 311790 560979 311824
rect 560945 311722 560979 311756
rect 561203 312606 561237 312640
rect 561203 312538 561237 312572
rect 561203 312470 561237 312504
rect 561203 312402 561237 312436
rect 561203 312334 561237 312368
rect 561203 312266 561237 312300
rect 561203 312198 561237 312232
rect 561203 312130 561237 312164
rect 561203 312062 561237 312096
rect 561203 311994 561237 312028
rect 561203 311926 561237 311960
rect 561203 311858 561237 311892
rect 561203 311790 561237 311824
rect 561203 311722 561237 311756
rect 561461 312606 561495 312640
rect 561461 312538 561495 312572
rect 561461 312470 561495 312504
rect 561461 312402 561495 312436
rect 561461 312334 561495 312368
rect 561461 312266 561495 312300
rect 561461 312198 561495 312232
rect 561461 312130 561495 312164
rect 561461 312062 561495 312096
rect 561461 311994 561495 312028
rect 561461 311926 561495 311960
rect 561461 311858 561495 311892
rect 561461 311790 561495 311824
rect 561461 311722 561495 311756
rect 561719 312606 561753 312640
rect 561719 312538 561753 312572
rect 561719 312470 561753 312504
rect 561719 312402 561753 312436
rect 561719 312334 561753 312368
rect 561719 312266 561753 312300
rect 561719 312198 561753 312232
rect 561719 312130 561753 312164
rect 561719 312062 561753 312096
rect 561719 311994 561753 312028
rect 561719 311926 561753 311960
rect 561719 311858 561753 311892
rect 561719 311790 561753 311824
rect 561719 311722 561753 311756
rect 561977 312606 562011 312640
rect 561977 312538 562011 312572
rect 561977 312470 562011 312504
rect 561977 312402 562011 312436
rect 561977 312334 562011 312368
rect 561977 312266 562011 312300
rect 561977 312198 562011 312232
rect 561977 312130 562011 312164
rect 561977 312062 562011 312096
rect 561977 311994 562011 312028
rect 561977 311926 562011 311960
rect 561977 311858 562011 311892
rect 561977 311790 562011 311824
rect 561977 311722 562011 311756
rect 562235 312606 562269 312640
rect 562235 312538 562269 312572
rect 562235 312470 562269 312504
rect 562235 312402 562269 312436
rect 562235 312334 562269 312368
rect 562235 312266 562269 312300
rect 562235 312198 562269 312232
rect 562235 312130 562269 312164
rect 562235 312062 562269 312096
rect 562235 311994 562269 312028
rect 562235 311926 562269 311960
rect 562235 311858 562269 311892
rect 562235 311790 562269 311824
rect 562235 311722 562269 311756
rect 562493 312606 562527 312640
rect 562493 312538 562527 312572
rect 562493 312470 562527 312504
rect 562493 312402 562527 312436
rect 562493 312334 562527 312368
rect 562493 312266 562527 312300
rect 562493 312198 562527 312232
rect 562493 312130 562527 312164
rect 562493 312062 562527 312096
rect 562493 311994 562527 312028
rect 562493 311926 562527 311960
rect 562493 311858 562527 311892
rect 562493 311790 562527 311824
rect 562493 311722 562527 311756
rect 562751 312606 562785 312640
rect 562751 312538 562785 312572
rect 562751 312470 562785 312504
rect 562751 312402 562785 312436
rect 562751 312334 562785 312368
rect 562751 312266 562785 312300
rect 562751 312198 562785 312232
rect 562751 312130 562785 312164
rect 562751 312062 562785 312096
rect 562751 311994 562785 312028
rect 562751 311926 562785 311960
rect 562751 311858 562785 311892
rect 562751 311790 562785 311824
rect 562751 311722 562785 311756
rect 563009 312606 563043 312640
rect 563009 312538 563043 312572
rect 563009 312470 563043 312504
rect 563009 312402 563043 312436
rect 563009 312334 563043 312368
rect 563009 312266 563043 312300
rect 563009 312198 563043 312232
rect 563009 312130 563043 312164
rect 563009 312062 563043 312096
rect 563009 311994 563043 312028
rect 563009 311926 563043 311960
rect 563009 311858 563043 311892
rect 563009 311790 563043 311824
rect 563009 311722 563043 311756
rect 563267 312606 563301 312640
rect 563267 312538 563301 312572
rect 563267 312470 563301 312504
rect 563267 312402 563301 312436
rect 563267 312334 563301 312368
rect 563267 312266 563301 312300
rect 563267 312198 563301 312232
rect 563267 312130 563301 312164
rect 563267 312062 563301 312096
rect 563267 311994 563301 312028
rect 563267 311926 563301 311960
rect 563267 311858 563301 311892
rect 563267 311790 563301 311824
rect 563267 311722 563301 311756
rect 563525 312606 563559 312640
rect 563525 312538 563559 312572
rect 563525 312470 563559 312504
rect 563525 312402 563559 312436
rect 563525 312334 563559 312368
rect 563525 312266 563559 312300
rect 563525 312198 563559 312232
rect 563525 312130 563559 312164
rect 563525 312062 563559 312096
rect 563525 311994 563559 312028
rect 563525 311926 563559 311960
rect 563525 311858 563559 311892
rect 563525 311790 563559 311824
rect 563525 311722 563559 311756
rect 563783 312606 563817 312640
rect 563783 312538 563817 312572
rect 563783 312470 563817 312504
rect 563783 312402 563817 312436
rect 563783 312334 563817 312368
rect 563783 312266 563817 312300
rect 563783 312198 563817 312232
rect 563783 312130 563817 312164
rect 563783 312062 563817 312096
rect 563783 311994 563817 312028
rect 563783 311926 563817 311960
rect 563783 311858 563817 311892
rect 563783 311790 563817 311824
rect 563783 311722 563817 311756
rect 564041 312606 564075 312640
rect 564041 312538 564075 312572
rect 564041 312470 564075 312504
rect 564041 312402 564075 312436
rect 564041 312334 564075 312368
rect 564041 312266 564075 312300
rect 564041 312198 564075 312232
rect 564041 312130 564075 312164
rect 564041 312062 564075 312096
rect 564041 311994 564075 312028
rect 564041 311926 564075 311960
rect 564041 311858 564075 311892
rect 564041 311790 564075 311824
rect 564041 311722 564075 311756
rect 564299 312606 564333 312640
rect 564299 312538 564333 312572
rect 564299 312470 564333 312504
rect 564299 312402 564333 312436
rect 564299 312334 564333 312368
rect 564299 312266 564333 312300
rect 564299 312198 564333 312232
rect 564299 312130 564333 312164
rect 564299 312062 564333 312096
rect 564299 311994 564333 312028
rect 564299 311926 564333 311960
rect 564299 311858 564333 311892
rect 564299 311790 564333 311824
rect 564299 311722 564333 311756
rect 564557 312606 564591 312640
rect 564557 312538 564591 312572
rect 564557 312470 564591 312504
rect 564557 312402 564591 312436
rect 564557 312334 564591 312368
rect 564557 312266 564591 312300
rect 564557 312198 564591 312232
rect 564557 312130 564591 312164
rect 564557 312062 564591 312096
rect 564557 311994 564591 312028
rect 564557 311926 564591 311960
rect 564557 311858 564591 311892
rect 564557 311790 564591 311824
rect 564557 311722 564591 311756
rect 564815 312606 564849 312640
rect 564815 312538 564849 312572
rect 564815 312470 564849 312504
rect 564815 312402 564849 312436
rect 564815 312334 564849 312368
rect 564815 312266 564849 312300
rect 564815 312198 564849 312232
rect 564815 312130 564849 312164
rect 564815 312062 564849 312096
rect 564815 311994 564849 312028
rect 564815 311926 564849 311960
rect 564815 311858 564849 311892
rect 564815 311790 564849 311824
rect 564815 311722 564849 311756
rect 565073 312606 565107 312640
rect 565073 312538 565107 312572
rect 565073 312470 565107 312504
rect 565073 312402 565107 312436
rect 565073 312334 565107 312368
rect 565073 312266 565107 312300
rect 565073 312198 565107 312232
rect 565073 312130 565107 312164
rect 565073 312062 565107 312096
rect 565073 311994 565107 312028
rect 565073 311926 565107 311960
rect 565073 311858 565107 311892
rect 565073 311790 565107 311824
rect 565073 311722 565107 311756
rect 565331 312606 565365 312640
rect 565331 312538 565365 312572
rect 565331 312470 565365 312504
rect 565331 312402 565365 312436
rect 565331 312334 565365 312368
rect 565331 312266 565365 312300
rect 565331 312198 565365 312232
rect 565331 312130 565365 312164
rect 565331 312062 565365 312096
rect 565331 311994 565365 312028
rect 565331 311926 565365 311960
rect 565331 311858 565365 311892
rect 565331 311790 565365 311824
rect 565331 311722 565365 311756
rect 565589 312606 565623 312640
rect 565589 312538 565623 312572
rect 565589 312470 565623 312504
rect 565589 312402 565623 312436
rect 565589 312334 565623 312368
rect 565589 312266 565623 312300
rect 565589 312198 565623 312232
rect 565589 312130 565623 312164
rect 565589 312062 565623 312096
rect 565589 311994 565623 312028
rect 565589 311926 565623 311960
rect 565589 311858 565623 311892
rect 565589 311790 565623 311824
rect 565589 311722 565623 311756
<< pdiffc >>
rect 575231 493148 575265 493182
rect 575231 493080 575265 493114
rect 575231 493012 575265 493046
rect 575231 492944 575265 492978
rect 575231 492876 575265 492910
rect 575231 492808 575265 492842
rect 575231 492740 575265 492774
rect 575231 492672 575265 492706
rect 575231 492604 575265 492638
rect 575231 492536 575265 492570
rect 575231 492468 575265 492502
rect 575231 492400 575265 492434
rect 575231 492332 575265 492366
rect 575231 492264 575265 492298
rect 575489 493148 575523 493182
rect 575489 493080 575523 493114
rect 575489 493012 575523 493046
rect 575489 492944 575523 492978
rect 575489 492876 575523 492910
rect 575489 492808 575523 492842
rect 575489 492740 575523 492774
rect 575489 492672 575523 492706
rect 575489 492604 575523 492638
rect 575489 492536 575523 492570
rect 575489 492468 575523 492502
rect 575489 492400 575523 492434
rect 575489 492332 575523 492366
rect 575489 492264 575523 492298
rect 575747 493148 575781 493182
rect 575747 493080 575781 493114
rect 575747 493012 575781 493046
rect 575747 492944 575781 492978
rect 575747 492876 575781 492910
rect 575747 492808 575781 492842
rect 575747 492740 575781 492774
rect 575747 492672 575781 492706
rect 575747 492604 575781 492638
rect 575747 492536 575781 492570
rect 575747 492468 575781 492502
rect 575747 492400 575781 492434
rect 575747 492332 575781 492366
rect 575747 492264 575781 492298
rect 576005 493148 576039 493182
rect 576005 493080 576039 493114
rect 576005 493012 576039 493046
rect 576005 492944 576039 492978
rect 576005 492876 576039 492910
rect 576005 492808 576039 492842
rect 576005 492740 576039 492774
rect 576005 492672 576039 492706
rect 576005 492604 576039 492638
rect 576005 492536 576039 492570
rect 576005 492468 576039 492502
rect 576005 492400 576039 492434
rect 576005 492332 576039 492366
rect 576005 492264 576039 492298
rect 576263 493148 576297 493182
rect 576263 493080 576297 493114
rect 576263 493012 576297 493046
rect 576263 492944 576297 492978
rect 576263 492876 576297 492910
rect 576263 492808 576297 492842
rect 576263 492740 576297 492774
rect 576263 492672 576297 492706
rect 576263 492604 576297 492638
rect 576263 492536 576297 492570
rect 576263 492468 576297 492502
rect 576263 492400 576297 492434
rect 576263 492332 576297 492366
rect 576263 492264 576297 492298
rect 576521 493148 576555 493182
rect 576521 493080 576555 493114
rect 576521 493012 576555 493046
rect 576521 492944 576555 492978
rect 576521 492876 576555 492910
rect 576521 492808 576555 492842
rect 576521 492740 576555 492774
rect 576521 492672 576555 492706
rect 576521 492604 576555 492638
rect 576521 492536 576555 492570
rect 576521 492468 576555 492502
rect 576521 492400 576555 492434
rect 576521 492332 576555 492366
rect 576521 492264 576555 492298
rect 576779 493148 576813 493182
rect 576779 493080 576813 493114
rect 576779 493012 576813 493046
rect 576779 492944 576813 492978
rect 576779 492876 576813 492910
rect 576779 492808 576813 492842
rect 576779 492740 576813 492774
rect 576779 492672 576813 492706
rect 576779 492604 576813 492638
rect 576779 492536 576813 492570
rect 576779 492468 576813 492502
rect 576779 492400 576813 492434
rect 576779 492332 576813 492366
rect 576779 492264 576813 492298
rect 577037 493148 577071 493182
rect 577037 493080 577071 493114
rect 577037 493012 577071 493046
rect 577037 492944 577071 492978
rect 577037 492876 577071 492910
rect 577037 492808 577071 492842
rect 577037 492740 577071 492774
rect 577037 492672 577071 492706
rect 577037 492604 577071 492638
rect 577037 492536 577071 492570
rect 577037 492468 577071 492502
rect 577037 492400 577071 492434
rect 577037 492332 577071 492366
rect 577037 492264 577071 492298
rect 577295 493148 577329 493182
rect 577295 493080 577329 493114
rect 577295 493012 577329 493046
rect 577295 492944 577329 492978
rect 577295 492876 577329 492910
rect 577295 492808 577329 492842
rect 577295 492740 577329 492774
rect 577295 492672 577329 492706
rect 577295 492604 577329 492638
rect 577295 492536 577329 492570
rect 577295 492468 577329 492502
rect 577295 492400 577329 492434
rect 577295 492332 577329 492366
rect 577295 492264 577329 492298
rect 577553 493148 577587 493182
rect 577553 493080 577587 493114
rect 577553 493012 577587 493046
rect 577553 492944 577587 492978
rect 577553 492876 577587 492910
rect 577553 492808 577587 492842
rect 577553 492740 577587 492774
rect 577553 492672 577587 492706
rect 577553 492604 577587 492638
rect 577553 492536 577587 492570
rect 577553 492468 577587 492502
rect 577553 492400 577587 492434
rect 577553 492332 577587 492366
rect 577553 492264 577587 492298
rect 577811 493148 577845 493182
rect 577811 493080 577845 493114
rect 577811 493012 577845 493046
rect 577811 492944 577845 492978
rect 577811 492876 577845 492910
rect 577811 492808 577845 492842
rect 577811 492740 577845 492774
rect 577811 492672 577845 492706
rect 577811 492604 577845 492638
rect 577811 492536 577845 492570
rect 577811 492468 577845 492502
rect 577811 492400 577845 492434
rect 577811 492332 577845 492366
rect 577811 492264 577845 492298
rect 578069 493148 578103 493182
rect 578069 493080 578103 493114
rect 578069 493012 578103 493046
rect 578069 492944 578103 492978
rect 578069 492876 578103 492910
rect 578069 492808 578103 492842
rect 578069 492740 578103 492774
rect 578069 492672 578103 492706
rect 578069 492604 578103 492638
rect 578069 492536 578103 492570
rect 578069 492468 578103 492502
rect 578069 492400 578103 492434
rect 578069 492332 578103 492366
rect 578069 492264 578103 492298
rect 578327 493148 578361 493182
rect 578327 493080 578361 493114
rect 578327 493012 578361 493046
rect 578327 492944 578361 492978
rect 578327 492876 578361 492910
rect 578327 492808 578361 492842
rect 578327 492740 578361 492774
rect 578327 492672 578361 492706
rect 578327 492604 578361 492638
rect 578327 492536 578361 492570
rect 578327 492468 578361 492502
rect 578327 492400 578361 492434
rect 578327 492332 578361 492366
rect 578327 492264 578361 492298
rect 578585 493148 578619 493182
rect 578585 493080 578619 493114
rect 578585 493012 578619 493046
rect 578585 492944 578619 492978
rect 578585 492876 578619 492910
rect 578585 492808 578619 492842
rect 578585 492740 578619 492774
rect 578585 492672 578619 492706
rect 578585 492604 578619 492638
rect 578585 492536 578619 492570
rect 578585 492468 578619 492502
rect 578585 492400 578619 492434
rect 578585 492332 578619 492366
rect 578585 492264 578619 492298
rect 578843 493148 578877 493182
rect 578843 493080 578877 493114
rect 578843 493012 578877 493046
rect 578843 492944 578877 492978
rect 578843 492876 578877 492910
rect 578843 492808 578877 492842
rect 578843 492740 578877 492774
rect 578843 492672 578877 492706
rect 578843 492604 578877 492638
rect 578843 492536 578877 492570
rect 578843 492468 578877 492502
rect 578843 492400 578877 492434
rect 578843 492332 578877 492366
rect 578843 492264 578877 492298
rect 579101 493148 579135 493182
rect 579101 493080 579135 493114
rect 579101 493012 579135 493046
rect 579101 492944 579135 492978
rect 579101 492876 579135 492910
rect 579101 492808 579135 492842
rect 579101 492740 579135 492774
rect 579101 492672 579135 492706
rect 579101 492604 579135 492638
rect 579101 492536 579135 492570
rect 579101 492468 579135 492502
rect 579101 492400 579135 492434
rect 579101 492332 579135 492366
rect 579101 492264 579135 492298
rect 579359 493148 579393 493182
rect 579359 493080 579393 493114
rect 579359 493012 579393 493046
rect 579359 492944 579393 492978
rect 579359 492876 579393 492910
rect 579359 492808 579393 492842
rect 579359 492740 579393 492774
rect 579359 492672 579393 492706
rect 579359 492604 579393 492638
rect 579359 492536 579393 492570
rect 579359 492468 579393 492502
rect 579359 492400 579393 492434
rect 579359 492332 579393 492366
rect 579359 492264 579393 492298
rect 579617 493148 579651 493182
rect 579617 493080 579651 493114
rect 579617 493012 579651 493046
rect 579617 492944 579651 492978
rect 579617 492876 579651 492910
rect 579617 492808 579651 492842
rect 579617 492740 579651 492774
rect 579617 492672 579651 492706
rect 579617 492604 579651 492638
rect 579617 492536 579651 492570
rect 579617 492468 579651 492502
rect 579617 492400 579651 492434
rect 579617 492332 579651 492366
rect 579617 492264 579651 492298
rect 579875 493148 579909 493182
rect 579875 493080 579909 493114
rect 579875 493012 579909 493046
rect 579875 492944 579909 492978
rect 579875 492876 579909 492910
rect 579875 492808 579909 492842
rect 579875 492740 579909 492774
rect 579875 492672 579909 492706
rect 579875 492604 579909 492638
rect 579875 492536 579909 492570
rect 579875 492468 579909 492502
rect 579875 492400 579909 492434
rect 579875 492332 579909 492366
rect 579875 492264 579909 492298
rect 580133 493148 580167 493182
rect 580133 493080 580167 493114
rect 580133 493012 580167 493046
rect 580133 492944 580167 492978
rect 580133 492876 580167 492910
rect 580133 492808 580167 492842
rect 580133 492740 580167 492774
rect 580133 492672 580167 492706
rect 580133 492604 580167 492638
rect 580133 492536 580167 492570
rect 580133 492468 580167 492502
rect 580133 492400 580167 492434
rect 580133 492332 580167 492366
rect 580133 492264 580167 492298
rect 580391 493148 580425 493182
rect 580391 493080 580425 493114
rect 580391 493012 580425 493046
rect 580391 492944 580425 492978
rect 580391 492876 580425 492910
rect 580391 492808 580425 492842
rect 580391 492740 580425 492774
rect 580391 492672 580425 492706
rect 580391 492604 580425 492638
rect 580391 492536 580425 492570
rect 580391 492468 580425 492502
rect 580391 492400 580425 492434
rect 580391 492332 580425 492366
rect 580391 492264 580425 492298
rect 574705 358844 574739 358878
rect 574705 358776 574739 358810
rect 574705 358708 574739 358742
rect 574705 358640 574739 358674
rect 574705 358572 574739 358606
rect 574705 358504 574739 358538
rect 574705 358436 574739 358470
rect 574705 358368 574739 358402
rect 574705 358300 574739 358334
rect 574705 358232 574739 358266
rect 574705 358164 574739 358198
rect 574705 358096 574739 358130
rect 574705 358028 574739 358062
rect 574705 357960 574739 357994
rect 574963 358844 574997 358878
rect 574963 358776 574997 358810
rect 574963 358708 574997 358742
rect 574963 358640 574997 358674
rect 574963 358572 574997 358606
rect 574963 358504 574997 358538
rect 574963 358436 574997 358470
rect 574963 358368 574997 358402
rect 574963 358300 574997 358334
rect 574963 358232 574997 358266
rect 574963 358164 574997 358198
rect 574963 358096 574997 358130
rect 574963 358028 574997 358062
rect 574963 357960 574997 357994
rect 575221 358844 575255 358878
rect 575221 358776 575255 358810
rect 575221 358708 575255 358742
rect 575221 358640 575255 358674
rect 575221 358572 575255 358606
rect 575221 358504 575255 358538
rect 575221 358436 575255 358470
rect 575221 358368 575255 358402
rect 575221 358300 575255 358334
rect 575221 358232 575255 358266
rect 575221 358164 575255 358198
rect 575221 358096 575255 358130
rect 575221 358028 575255 358062
rect 575221 357960 575255 357994
rect 575479 358844 575513 358878
rect 575479 358776 575513 358810
rect 575479 358708 575513 358742
rect 575479 358640 575513 358674
rect 575479 358572 575513 358606
rect 575479 358504 575513 358538
rect 575479 358436 575513 358470
rect 575479 358368 575513 358402
rect 575479 358300 575513 358334
rect 575479 358232 575513 358266
rect 575479 358164 575513 358198
rect 575479 358096 575513 358130
rect 575479 358028 575513 358062
rect 575479 357960 575513 357994
rect 575737 358844 575771 358878
rect 575737 358776 575771 358810
rect 575737 358708 575771 358742
rect 575737 358640 575771 358674
rect 575737 358572 575771 358606
rect 575737 358504 575771 358538
rect 575737 358436 575771 358470
rect 575737 358368 575771 358402
rect 575737 358300 575771 358334
rect 575737 358232 575771 358266
rect 575737 358164 575771 358198
rect 575737 358096 575771 358130
rect 575737 358028 575771 358062
rect 575737 357960 575771 357994
rect 575995 358844 576029 358878
rect 575995 358776 576029 358810
rect 575995 358708 576029 358742
rect 575995 358640 576029 358674
rect 575995 358572 576029 358606
rect 575995 358504 576029 358538
rect 575995 358436 576029 358470
rect 575995 358368 576029 358402
rect 575995 358300 576029 358334
rect 575995 358232 576029 358266
rect 575995 358164 576029 358198
rect 575995 358096 576029 358130
rect 575995 358028 576029 358062
rect 575995 357960 576029 357994
rect 576253 358844 576287 358878
rect 576253 358776 576287 358810
rect 576253 358708 576287 358742
rect 576253 358640 576287 358674
rect 576253 358572 576287 358606
rect 576253 358504 576287 358538
rect 576253 358436 576287 358470
rect 576253 358368 576287 358402
rect 576253 358300 576287 358334
rect 576253 358232 576287 358266
rect 576253 358164 576287 358198
rect 576253 358096 576287 358130
rect 576253 358028 576287 358062
rect 576253 357960 576287 357994
rect 576511 358844 576545 358878
rect 576511 358776 576545 358810
rect 576511 358708 576545 358742
rect 576511 358640 576545 358674
rect 576511 358572 576545 358606
rect 576511 358504 576545 358538
rect 576511 358436 576545 358470
rect 576511 358368 576545 358402
rect 576511 358300 576545 358334
rect 576511 358232 576545 358266
rect 576511 358164 576545 358198
rect 576511 358096 576545 358130
rect 576511 358028 576545 358062
rect 576511 357960 576545 357994
rect 576769 358844 576803 358878
rect 576769 358776 576803 358810
rect 576769 358708 576803 358742
rect 576769 358640 576803 358674
rect 576769 358572 576803 358606
rect 576769 358504 576803 358538
rect 576769 358436 576803 358470
rect 576769 358368 576803 358402
rect 576769 358300 576803 358334
rect 576769 358232 576803 358266
rect 576769 358164 576803 358198
rect 576769 358096 576803 358130
rect 576769 358028 576803 358062
rect 576769 357960 576803 357994
rect 577027 358844 577061 358878
rect 577027 358776 577061 358810
rect 577027 358708 577061 358742
rect 577027 358640 577061 358674
rect 577027 358572 577061 358606
rect 577027 358504 577061 358538
rect 577027 358436 577061 358470
rect 577027 358368 577061 358402
rect 577027 358300 577061 358334
rect 577027 358232 577061 358266
rect 577027 358164 577061 358198
rect 577027 358096 577061 358130
rect 577027 358028 577061 358062
rect 577027 357960 577061 357994
rect 577285 358844 577319 358878
rect 577285 358776 577319 358810
rect 577285 358708 577319 358742
rect 577285 358640 577319 358674
rect 577285 358572 577319 358606
rect 577285 358504 577319 358538
rect 577285 358436 577319 358470
rect 577285 358368 577319 358402
rect 577285 358300 577319 358334
rect 577285 358232 577319 358266
rect 577285 358164 577319 358198
rect 577285 358096 577319 358130
rect 577285 358028 577319 358062
rect 577285 357960 577319 357994
rect 577543 358844 577577 358878
rect 577543 358776 577577 358810
rect 577543 358708 577577 358742
rect 577543 358640 577577 358674
rect 577543 358572 577577 358606
rect 577543 358504 577577 358538
rect 577543 358436 577577 358470
rect 577543 358368 577577 358402
rect 577543 358300 577577 358334
rect 577543 358232 577577 358266
rect 577543 358164 577577 358198
rect 577543 358096 577577 358130
rect 577543 358028 577577 358062
rect 577543 357960 577577 357994
rect 577801 358844 577835 358878
rect 577801 358776 577835 358810
rect 577801 358708 577835 358742
rect 577801 358640 577835 358674
rect 577801 358572 577835 358606
rect 577801 358504 577835 358538
rect 577801 358436 577835 358470
rect 577801 358368 577835 358402
rect 577801 358300 577835 358334
rect 577801 358232 577835 358266
rect 577801 358164 577835 358198
rect 577801 358096 577835 358130
rect 577801 358028 577835 358062
rect 577801 357960 577835 357994
rect 578059 358844 578093 358878
rect 578059 358776 578093 358810
rect 578059 358708 578093 358742
rect 578059 358640 578093 358674
rect 578059 358572 578093 358606
rect 578059 358504 578093 358538
rect 578059 358436 578093 358470
rect 578059 358368 578093 358402
rect 578059 358300 578093 358334
rect 578059 358232 578093 358266
rect 578059 358164 578093 358198
rect 578059 358096 578093 358130
rect 578059 358028 578093 358062
rect 578059 357960 578093 357994
rect 578317 358844 578351 358878
rect 578317 358776 578351 358810
rect 578317 358708 578351 358742
rect 578317 358640 578351 358674
rect 578317 358572 578351 358606
rect 578317 358504 578351 358538
rect 578317 358436 578351 358470
rect 578317 358368 578351 358402
rect 578317 358300 578351 358334
rect 578317 358232 578351 358266
rect 578317 358164 578351 358198
rect 578317 358096 578351 358130
rect 578317 358028 578351 358062
rect 578317 357960 578351 357994
rect 578575 358844 578609 358878
rect 578575 358776 578609 358810
rect 578575 358708 578609 358742
rect 578575 358640 578609 358674
rect 578575 358572 578609 358606
rect 578575 358504 578609 358538
rect 578575 358436 578609 358470
rect 578575 358368 578609 358402
rect 578575 358300 578609 358334
rect 578575 358232 578609 358266
rect 578575 358164 578609 358198
rect 578575 358096 578609 358130
rect 578575 358028 578609 358062
rect 578575 357960 578609 357994
rect 578833 358844 578867 358878
rect 578833 358776 578867 358810
rect 578833 358708 578867 358742
rect 578833 358640 578867 358674
rect 578833 358572 578867 358606
rect 578833 358504 578867 358538
rect 578833 358436 578867 358470
rect 578833 358368 578867 358402
rect 578833 358300 578867 358334
rect 578833 358232 578867 358266
rect 578833 358164 578867 358198
rect 578833 358096 578867 358130
rect 578833 358028 578867 358062
rect 578833 357960 578867 357994
rect 579091 358844 579125 358878
rect 579091 358776 579125 358810
rect 579091 358708 579125 358742
rect 579091 358640 579125 358674
rect 579091 358572 579125 358606
rect 579091 358504 579125 358538
rect 579091 358436 579125 358470
rect 579091 358368 579125 358402
rect 579091 358300 579125 358334
rect 579091 358232 579125 358266
rect 579091 358164 579125 358198
rect 579091 358096 579125 358130
rect 579091 358028 579125 358062
rect 579091 357960 579125 357994
rect 579349 358844 579383 358878
rect 579349 358776 579383 358810
rect 579349 358708 579383 358742
rect 579349 358640 579383 358674
rect 579349 358572 579383 358606
rect 579349 358504 579383 358538
rect 579349 358436 579383 358470
rect 579349 358368 579383 358402
rect 579349 358300 579383 358334
rect 579349 358232 579383 358266
rect 579349 358164 579383 358198
rect 579349 358096 579383 358130
rect 579349 358028 579383 358062
rect 579349 357960 579383 357994
rect 579607 358844 579641 358878
rect 579607 358776 579641 358810
rect 579607 358708 579641 358742
rect 579607 358640 579641 358674
rect 579607 358572 579641 358606
rect 579607 358504 579641 358538
rect 579607 358436 579641 358470
rect 579607 358368 579641 358402
rect 579607 358300 579641 358334
rect 579607 358232 579641 358266
rect 579607 358164 579641 358198
rect 579607 358096 579641 358130
rect 579607 358028 579641 358062
rect 579607 357960 579641 357994
rect 579865 358844 579899 358878
rect 579865 358776 579899 358810
rect 579865 358708 579899 358742
rect 579865 358640 579899 358674
rect 579865 358572 579899 358606
rect 579865 358504 579899 358538
rect 579865 358436 579899 358470
rect 579865 358368 579899 358402
rect 579865 358300 579899 358334
rect 579865 358232 579899 358266
rect 579865 358164 579899 358198
rect 579865 358096 579899 358130
rect 579865 358028 579899 358062
rect 579865 357960 579899 357994
rect 575153 312676 575187 312710
rect 575153 312608 575187 312642
rect 575153 312540 575187 312574
rect 575153 312472 575187 312506
rect 575153 312404 575187 312438
rect 575153 312336 575187 312370
rect 575153 312268 575187 312302
rect 575153 312200 575187 312234
rect 575153 312132 575187 312166
rect 575153 312064 575187 312098
rect 575153 311996 575187 312030
rect 575153 311928 575187 311962
rect 575153 311860 575187 311894
rect 575153 311792 575187 311826
rect 575411 312676 575445 312710
rect 575411 312608 575445 312642
rect 575411 312540 575445 312574
rect 575411 312472 575445 312506
rect 575411 312404 575445 312438
rect 575411 312336 575445 312370
rect 575411 312268 575445 312302
rect 575411 312200 575445 312234
rect 575411 312132 575445 312166
rect 575411 312064 575445 312098
rect 575411 311996 575445 312030
rect 575411 311928 575445 311962
rect 575411 311860 575445 311894
rect 575411 311792 575445 311826
rect 575669 312676 575703 312710
rect 575669 312608 575703 312642
rect 575669 312540 575703 312574
rect 575669 312472 575703 312506
rect 575669 312404 575703 312438
rect 575669 312336 575703 312370
rect 575669 312268 575703 312302
rect 575669 312200 575703 312234
rect 575669 312132 575703 312166
rect 575669 312064 575703 312098
rect 575669 311996 575703 312030
rect 575669 311928 575703 311962
rect 575669 311860 575703 311894
rect 575669 311792 575703 311826
rect 575927 312676 575961 312710
rect 575927 312608 575961 312642
rect 575927 312540 575961 312574
rect 575927 312472 575961 312506
rect 575927 312404 575961 312438
rect 575927 312336 575961 312370
rect 575927 312268 575961 312302
rect 575927 312200 575961 312234
rect 575927 312132 575961 312166
rect 575927 312064 575961 312098
rect 575927 311996 575961 312030
rect 575927 311928 575961 311962
rect 575927 311860 575961 311894
rect 575927 311792 575961 311826
rect 576185 312676 576219 312710
rect 576185 312608 576219 312642
rect 576185 312540 576219 312574
rect 576185 312472 576219 312506
rect 576185 312404 576219 312438
rect 576185 312336 576219 312370
rect 576185 312268 576219 312302
rect 576185 312200 576219 312234
rect 576185 312132 576219 312166
rect 576185 312064 576219 312098
rect 576185 311996 576219 312030
rect 576185 311928 576219 311962
rect 576185 311860 576219 311894
rect 576185 311792 576219 311826
rect 576443 312676 576477 312710
rect 576443 312608 576477 312642
rect 576443 312540 576477 312574
rect 576443 312472 576477 312506
rect 576443 312404 576477 312438
rect 576443 312336 576477 312370
rect 576443 312268 576477 312302
rect 576443 312200 576477 312234
rect 576443 312132 576477 312166
rect 576443 312064 576477 312098
rect 576443 311996 576477 312030
rect 576443 311928 576477 311962
rect 576443 311860 576477 311894
rect 576443 311792 576477 311826
rect 576701 312676 576735 312710
rect 576701 312608 576735 312642
rect 576701 312540 576735 312574
rect 576701 312472 576735 312506
rect 576701 312404 576735 312438
rect 576701 312336 576735 312370
rect 576701 312268 576735 312302
rect 576701 312200 576735 312234
rect 576701 312132 576735 312166
rect 576701 312064 576735 312098
rect 576701 311996 576735 312030
rect 576701 311928 576735 311962
rect 576701 311860 576735 311894
rect 576701 311792 576735 311826
rect 576959 312676 576993 312710
rect 576959 312608 576993 312642
rect 576959 312540 576993 312574
rect 576959 312472 576993 312506
rect 576959 312404 576993 312438
rect 576959 312336 576993 312370
rect 576959 312268 576993 312302
rect 576959 312200 576993 312234
rect 576959 312132 576993 312166
rect 576959 312064 576993 312098
rect 576959 311996 576993 312030
rect 576959 311928 576993 311962
rect 576959 311860 576993 311894
rect 576959 311792 576993 311826
rect 577217 312676 577251 312710
rect 577217 312608 577251 312642
rect 577217 312540 577251 312574
rect 577217 312472 577251 312506
rect 577217 312404 577251 312438
rect 577217 312336 577251 312370
rect 577217 312268 577251 312302
rect 577217 312200 577251 312234
rect 577217 312132 577251 312166
rect 577217 312064 577251 312098
rect 577217 311996 577251 312030
rect 577217 311928 577251 311962
rect 577217 311860 577251 311894
rect 577217 311792 577251 311826
rect 577475 312676 577509 312710
rect 577475 312608 577509 312642
rect 577475 312540 577509 312574
rect 577475 312472 577509 312506
rect 577475 312404 577509 312438
rect 577475 312336 577509 312370
rect 577475 312268 577509 312302
rect 577475 312200 577509 312234
rect 577475 312132 577509 312166
rect 577475 312064 577509 312098
rect 577475 311996 577509 312030
rect 577475 311928 577509 311962
rect 577475 311860 577509 311894
rect 577475 311792 577509 311826
rect 577733 312676 577767 312710
rect 577733 312608 577767 312642
rect 577733 312540 577767 312574
rect 577733 312472 577767 312506
rect 577733 312404 577767 312438
rect 577733 312336 577767 312370
rect 577733 312268 577767 312302
rect 577733 312200 577767 312234
rect 577733 312132 577767 312166
rect 577733 312064 577767 312098
rect 577733 311996 577767 312030
rect 577733 311928 577767 311962
rect 577733 311860 577767 311894
rect 577733 311792 577767 311826
rect 577991 312676 578025 312710
rect 577991 312608 578025 312642
rect 577991 312540 578025 312574
rect 577991 312472 578025 312506
rect 577991 312404 578025 312438
rect 577991 312336 578025 312370
rect 577991 312268 578025 312302
rect 577991 312200 578025 312234
rect 577991 312132 578025 312166
rect 577991 312064 578025 312098
rect 577991 311996 578025 312030
rect 577991 311928 578025 311962
rect 577991 311860 578025 311894
rect 577991 311792 578025 311826
rect 578249 312676 578283 312710
rect 578249 312608 578283 312642
rect 578249 312540 578283 312574
rect 578249 312472 578283 312506
rect 578249 312404 578283 312438
rect 578249 312336 578283 312370
rect 578249 312268 578283 312302
rect 578249 312200 578283 312234
rect 578249 312132 578283 312166
rect 578249 312064 578283 312098
rect 578249 311996 578283 312030
rect 578249 311928 578283 311962
rect 578249 311860 578283 311894
rect 578249 311792 578283 311826
rect 578507 312676 578541 312710
rect 578507 312608 578541 312642
rect 578507 312540 578541 312574
rect 578507 312472 578541 312506
rect 578507 312404 578541 312438
rect 578507 312336 578541 312370
rect 578507 312268 578541 312302
rect 578507 312200 578541 312234
rect 578507 312132 578541 312166
rect 578507 312064 578541 312098
rect 578507 311996 578541 312030
rect 578507 311928 578541 311962
rect 578507 311860 578541 311894
rect 578507 311792 578541 311826
rect 578765 312676 578799 312710
rect 578765 312608 578799 312642
rect 578765 312540 578799 312574
rect 578765 312472 578799 312506
rect 578765 312404 578799 312438
rect 578765 312336 578799 312370
rect 578765 312268 578799 312302
rect 578765 312200 578799 312234
rect 578765 312132 578799 312166
rect 578765 312064 578799 312098
rect 578765 311996 578799 312030
rect 578765 311928 578799 311962
rect 578765 311860 578799 311894
rect 578765 311792 578799 311826
rect 579023 312676 579057 312710
rect 579023 312608 579057 312642
rect 579023 312540 579057 312574
rect 579023 312472 579057 312506
rect 579023 312404 579057 312438
rect 579023 312336 579057 312370
rect 579023 312268 579057 312302
rect 579023 312200 579057 312234
rect 579023 312132 579057 312166
rect 579023 312064 579057 312098
rect 579023 311996 579057 312030
rect 579023 311928 579057 311962
rect 579023 311860 579057 311894
rect 579023 311792 579057 311826
rect 579281 312676 579315 312710
rect 579281 312608 579315 312642
rect 579281 312540 579315 312574
rect 579281 312472 579315 312506
rect 579281 312404 579315 312438
rect 579281 312336 579315 312370
rect 579281 312268 579315 312302
rect 579281 312200 579315 312234
rect 579281 312132 579315 312166
rect 579281 312064 579315 312098
rect 579281 311996 579315 312030
rect 579281 311928 579315 311962
rect 579281 311860 579315 311894
rect 579281 311792 579315 311826
rect 579539 312676 579573 312710
rect 579539 312608 579573 312642
rect 579539 312540 579573 312574
rect 579539 312472 579573 312506
rect 579539 312404 579573 312438
rect 579539 312336 579573 312370
rect 579539 312268 579573 312302
rect 579539 312200 579573 312234
rect 579539 312132 579573 312166
rect 579539 312064 579573 312098
rect 579539 311996 579573 312030
rect 579539 311928 579573 311962
rect 579539 311860 579573 311894
rect 579539 311792 579573 311826
rect 579797 312676 579831 312710
rect 579797 312608 579831 312642
rect 579797 312540 579831 312574
rect 579797 312472 579831 312506
rect 579797 312404 579831 312438
rect 579797 312336 579831 312370
rect 579797 312268 579831 312302
rect 579797 312200 579831 312234
rect 579797 312132 579831 312166
rect 579797 312064 579831 312098
rect 579797 311996 579831 312030
rect 579797 311928 579831 311962
rect 579797 311860 579831 311894
rect 579797 311792 579831 311826
rect 580055 312676 580089 312710
rect 580055 312608 580089 312642
rect 580055 312540 580089 312574
rect 580055 312472 580089 312506
rect 580055 312404 580089 312438
rect 580055 312336 580089 312370
rect 580055 312268 580089 312302
rect 580055 312200 580089 312234
rect 580055 312132 580089 312166
rect 580055 312064 580089 312098
rect 580055 311996 580089 312030
rect 580055 311928 580089 311962
rect 580055 311860 580089 311894
rect 580055 311792 580089 311826
rect 580313 312676 580347 312710
rect 580313 312608 580347 312642
rect 580313 312540 580347 312574
rect 580313 312472 580347 312506
rect 580313 312404 580347 312438
rect 580313 312336 580347 312370
rect 580313 312268 580347 312302
rect 580313 312200 580347 312234
rect 580313 312132 580347 312166
rect 580313 312064 580347 312098
rect 580313 311996 580347 312030
rect 580313 311928 580347 311962
rect 580313 311860 580347 311894
rect 580313 311792 580347 311826
<< psubdiff >>
rect 565900 492106 565940 492149
rect 562162 492076 562282 492079
rect 562162 492042 562203 492076
rect 562237 492042 562282 492076
rect 562162 492029 562282 492042
rect 563462 492076 563582 492079
rect 563462 492042 563503 492076
rect 563537 492042 563582 492076
rect 563462 492029 563582 492042
rect 564762 492076 564882 492079
rect 564762 492042 564803 492076
rect 564837 492042 564882 492076
rect 564762 492029 564882 492042
rect 565900 492072 565903 492106
rect 565937 492072 565940 492106
rect 565900 492029 565940 492072
rect 565836 402964 565876 403007
rect 562098 402934 562218 402937
rect 562098 402900 562139 402934
rect 562173 402900 562218 402934
rect 562098 402887 562218 402900
rect 563398 402934 563518 402937
rect 563398 402900 563439 402934
rect 563473 402900 563518 402934
rect 563398 402887 563518 402900
rect 564698 402934 564818 402937
rect 564698 402900 564739 402934
rect 564773 402900 564818 402934
rect 564698 402887 564818 402900
rect 565836 402930 565839 402964
rect 565873 402930 565876 402964
rect 565836 402887 565876 402930
rect 565792 357646 565832 357689
rect 562054 357616 562174 357619
rect 562054 357582 562095 357616
rect 562129 357582 562174 357616
rect 562054 357569 562174 357582
rect 563354 357616 563474 357619
rect 563354 357582 563395 357616
rect 563429 357582 563474 357616
rect 563354 357569 563474 357582
rect 564654 357616 564774 357619
rect 564654 357582 564695 357616
rect 564729 357582 564774 357616
rect 564654 357569 564774 357582
rect 565792 357612 565795 357646
rect 565829 357612 565832 357646
rect 565792 357569 565832 357612
rect 565654 311338 565694 311381
rect 561916 311308 562036 311311
rect 561916 311274 561957 311308
rect 561991 311274 562036 311308
rect 561916 311261 562036 311274
rect 563216 311308 563336 311311
rect 563216 311274 563257 311308
rect 563291 311274 563336 311308
rect 563216 311261 563336 311274
rect 564516 311308 564636 311311
rect 564516 311274 564557 311308
rect 564591 311274 564636 311308
rect 564516 311261 564636 311274
rect 565654 311304 565657 311338
rect 565691 311304 565694 311338
rect 565654 311261 565694 311304
<< nsubdiff >>
rect 576754 493530 576874 493533
rect 576754 493496 576795 493530
rect 576829 493496 576874 493530
rect 576754 493493 576874 493496
rect 578054 493530 578174 493533
rect 578054 493496 578095 493530
rect 578129 493496 578174 493530
rect 578054 493493 578174 493496
rect 579354 493530 579474 493533
rect 579354 493496 579395 493530
rect 579429 493496 579474 493530
rect 579354 493493 579474 493496
rect 580492 493480 580532 493523
rect 580492 493446 580495 493480
rect 580529 493446 580532 493480
rect 580492 493403 580532 493446
rect 576228 359226 576348 359229
rect 576228 359192 576269 359226
rect 576303 359192 576348 359226
rect 576228 359189 576348 359192
rect 577528 359226 577648 359229
rect 577528 359192 577569 359226
rect 577603 359192 577648 359226
rect 577528 359189 577648 359192
rect 578828 359226 578948 359229
rect 578828 359192 578869 359226
rect 578903 359192 578948 359226
rect 578828 359189 578948 359192
rect 579966 359176 580006 359219
rect 579966 359142 579969 359176
rect 580003 359142 580006 359176
rect 579966 359099 580006 359142
rect 576676 313058 576796 313061
rect 576676 313024 576717 313058
rect 576751 313024 576796 313058
rect 576676 313021 576796 313024
rect 577976 313058 578096 313061
rect 577976 313024 578017 313058
rect 578051 313024 578096 313058
rect 577976 313021 578096 313024
rect 579276 313058 579396 313061
rect 579276 313024 579317 313058
rect 579351 313024 579396 313058
rect 579276 313021 579396 313024
rect 580414 313008 580454 313051
rect 580414 312974 580417 313008
rect 580451 312974 580454 313008
rect 580414 312931 580454 312974
<< psubdiffcont >>
rect 562203 492042 562237 492076
rect 563503 492042 563537 492076
rect 564803 492042 564837 492076
rect 565903 492072 565937 492106
rect 562139 402900 562173 402934
rect 563439 402900 563473 402934
rect 564739 402900 564773 402934
rect 565839 402930 565873 402964
rect 562095 357582 562129 357616
rect 563395 357582 563429 357616
rect 564695 357582 564729 357616
rect 565795 357612 565829 357646
rect 561957 311274 561991 311308
rect 563257 311274 563291 311308
rect 564557 311274 564591 311308
rect 565657 311304 565691 311338
<< nsubdiffcont >>
rect 576795 493496 576829 493530
rect 578095 493496 578129 493530
rect 579395 493496 579429 493530
rect 580495 493446 580529 493480
rect 576269 359192 576303 359226
rect 577569 359192 577603 359226
rect 578869 359192 578903 359226
rect 579969 359142 580003 359176
rect 576717 313024 576751 313058
rect 578017 313024 578051 313058
rect 579317 313024 579351 313058
rect 580417 312974 580451 313008
<< poly >>
rect 560721 493449 560921 493475
rect 560979 493449 561179 493475
rect 561237 493449 561437 493475
rect 561495 493449 561695 493475
rect 561753 493449 561953 493475
rect 562011 493449 562211 493475
rect 562269 493449 562469 493475
rect 562527 493449 562727 493475
rect 562785 493449 562985 493475
rect 563043 493449 563243 493475
rect 563301 493449 563501 493475
rect 563559 493449 563759 493475
rect 563817 493449 564017 493475
rect 564075 493449 564275 493475
rect 564333 493449 564533 493475
rect 564591 493449 564791 493475
rect 564849 493449 565049 493475
rect 565107 493449 565307 493475
rect 565365 493449 565565 493475
rect 565623 493449 565823 493475
rect 575277 493223 575477 493249
rect 575535 493223 575735 493249
rect 575793 493223 575993 493249
rect 576051 493223 576251 493249
rect 576309 493223 576509 493249
rect 576567 493223 576767 493249
rect 576825 493223 577025 493249
rect 577083 493223 577283 493249
rect 577341 493223 577541 493249
rect 577599 493223 577799 493249
rect 577857 493223 578057 493249
rect 578115 493223 578315 493249
rect 578373 493223 578573 493249
rect 578631 493223 578831 493249
rect 578889 493223 579089 493249
rect 579147 493223 579347 493249
rect 579405 493223 579605 493249
rect 579663 493223 579863 493249
rect 579921 493223 580121 493249
rect 580179 493223 580379 493249
rect 560721 492423 560921 492449
rect 560979 492423 561179 492449
rect 561237 492423 561437 492449
rect 561495 492423 561695 492449
rect 561753 492423 561953 492449
rect 562011 492423 562211 492449
rect 562269 492423 562469 492449
rect 562527 492423 562727 492449
rect 562785 492423 562985 492449
rect 563043 492423 563243 492449
rect 563301 492423 563501 492449
rect 563559 492423 563759 492449
rect 563817 492423 564017 492449
rect 564075 492423 564275 492449
rect 564333 492423 564533 492449
rect 564591 492423 564791 492449
rect 564849 492423 565049 492449
rect 565107 492423 565307 492449
rect 565365 492423 565565 492449
rect 565623 492423 565823 492449
rect 560776 492233 560896 492423
rect 561032 492233 561152 492423
rect 561288 492233 561408 492423
rect 561544 492233 561664 492423
rect 561800 492233 561920 492423
rect 562056 492233 562176 492423
rect 562312 492233 562432 492423
rect 562568 492233 562688 492423
rect 562824 492233 562944 492423
rect 563080 492233 563200 492423
rect 563336 492233 563456 492423
rect 563592 492233 563712 492423
rect 563848 492233 563968 492423
rect 564104 492233 564224 492423
rect 564360 492233 564480 492423
rect 564616 492233 564736 492423
rect 564872 492233 564992 492423
rect 565128 492233 565248 492423
rect 565384 492233 565504 492423
rect 565640 492233 565760 492423
rect 560664 492200 565800 492233
rect 560664 492166 560863 492200
rect 560897 492166 561063 492200
rect 561097 492166 561263 492200
rect 561297 492166 561463 492200
rect 561497 492166 561663 492200
rect 561697 492166 561863 492200
rect 561897 492166 562063 492200
rect 562097 492166 562263 492200
rect 562297 492166 562463 492200
rect 562497 492166 562663 492200
rect 562697 492166 562863 492200
rect 562897 492166 563063 492200
rect 563097 492166 563263 492200
rect 563297 492166 563463 492200
rect 563497 492166 563663 492200
rect 563697 492166 563863 492200
rect 563897 492166 564063 492200
rect 564097 492166 564263 492200
rect 564297 492166 564463 492200
rect 564497 492166 564663 492200
rect 564697 492166 564863 492200
rect 564897 492166 565063 492200
rect 565097 492166 565263 492200
rect 565297 492166 565463 492200
rect 565497 492166 565663 492200
rect 565697 492166 565800 492200
rect 575277 492197 575477 492223
rect 575535 492197 575735 492223
rect 575793 492197 575993 492223
rect 576051 492197 576251 492223
rect 576309 492197 576509 492223
rect 576567 492197 576767 492223
rect 576825 492197 577025 492223
rect 577083 492197 577283 492223
rect 577341 492197 577541 492223
rect 577599 492197 577799 492223
rect 577857 492197 578057 492223
rect 578115 492197 578315 492223
rect 578373 492197 578573 492223
rect 578631 492197 578831 492223
rect 578889 492197 579089 492223
rect 579147 492197 579347 492223
rect 579405 492197 579605 492223
rect 579663 492197 579863 492223
rect 579921 492197 580121 492223
rect 580179 492197 580379 492223
rect 560664 492133 565800 492166
rect 575348 491951 575468 492197
rect 575604 491951 575724 492197
rect 575860 491951 575980 492197
rect 576116 491951 576236 492197
rect 576372 491951 576492 492197
rect 576628 491951 576748 492197
rect 576884 491951 577004 492197
rect 577140 491951 577260 492197
rect 577396 491951 577516 492197
rect 577652 491951 577772 492197
rect 577908 491951 578028 492197
rect 578164 491951 578284 492197
rect 578420 491951 578540 492197
rect 578676 491951 578796 492197
rect 578932 491951 579052 492197
rect 579188 491951 579308 492197
rect 579444 491951 579564 492197
rect 579700 491951 579820 492197
rect 579956 491951 580076 492197
rect 580212 491951 580332 492197
rect 575184 491918 580472 491951
rect 575184 491884 575255 491918
rect 575289 491884 575455 491918
rect 575489 491884 575655 491918
rect 575689 491884 575855 491918
rect 575889 491884 576055 491918
rect 576089 491884 576255 491918
rect 576289 491884 576455 491918
rect 576489 491884 576655 491918
rect 576689 491884 576855 491918
rect 576889 491884 577055 491918
rect 577089 491884 577255 491918
rect 577289 491884 577455 491918
rect 577489 491884 577655 491918
rect 577689 491884 577855 491918
rect 577889 491884 578055 491918
rect 578089 491884 578255 491918
rect 578289 491884 578455 491918
rect 578489 491884 578655 491918
rect 578689 491884 578855 491918
rect 578889 491884 579055 491918
rect 579089 491884 579255 491918
rect 579289 491884 579455 491918
rect 579489 491884 579655 491918
rect 579689 491884 579855 491918
rect 579889 491884 580055 491918
rect 580089 491884 580255 491918
rect 580289 491884 580472 491918
rect 575184 491851 580472 491884
rect 560657 404307 560857 404333
rect 560915 404307 561115 404333
rect 561173 404307 561373 404333
rect 561431 404307 561631 404333
rect 561689 404307 561889 404333
rect 561947 404307 562147 404333
rect 562205 404307 562405 404333
rect 562463 404307 562663 404333
rect 562721 404307 562921 404333
rect 562979 404307 563179 404333
rect 563237 404307 563437 404333
rect 563495 404307 563695 404333
rect 563753 404307 563953 404333
rect 564011 404307 564211 404333
rect 564269 404307 564469 404333
rect 564527 404307 564727 404333
rect 564785 404307 564985 404333
rect 565043 404307 565243 404333
rect 565301 404307 565501 404333
rect 565559 404307 565759 404333
rect 560657 403281 560857 403307
rect 560915 403281 561115 403307
rect 561173 403281 561373 403307
rect 561431 403281 561631 403307
rect 561689 403281 561889 403307
rect 561947 403281 562147 403307
rect 562205 403281 562405 403307
rect 562463 403281 562663 403307
rect 562721 403281 562921 403307
rect 562979 403281 563179 403307
rect 563237 403281 563437 403307
rect 563495 403281 563695 403307
rect 563753 403281 563953 403307
rect 564011 403281 564211 403307
rect 564269 403281 564469 403307
rect 564527 403281 564727 403307
rect 564785 403281 564985 403307
rect 565043 403281 565243 403307
rect 565301 403281 565501 403307
rect 565559 403281 565759 403307
rect 560712 403091 560832 403281
rect 560968 403091 561088 403281
rect 561224 403091 561344 403281
rect 561480 403091 561600 403281
rect 561736 403091 561856 403281
rect 561992 403091 562112 403281
rect 562248 403091 562368 403281
rect 562504 403091 562624 403281
rect 562760 403091 562880 403281
rect 563016 403091 563136 403281
rect 563272 403091 563392 403281
rect 563528 403091 563648 403281
rect 563784 403091 563904 403281
rect 564040 403091 564160 403281
rect 564296 403091 564416 403281
rect 564552 403091 564672 403281
rect 564808 403091 564928 403281
rect 565064 403091 565184 403281
rect 565320 403091 565440 403281
rect 565576 403091 565696 403281
rect 560600 403058 565736 403091
rect 560600 403024 560799 403058
rect 560833 403024 560999 403058
rect 561033 403024 561199 403058
rect 561233 403024 561399 403058
rect 561433 403024 561599 403058
rect 561633 403024 561799 403058
rect 561833 403024 561999 403058
rect 562033 403024 562199 403058
rect 562233 403024 562399 403058
rect 562433 403024 562599 403058
rect 562633 403024 562799 403058
rect 562833 403024 562999 403058
rect 563033 403024 563199 403058
rect 563233 403024 563399 403058
rect 563433 403024 563599 403058
rect 563633 403024 563799 403058
rect 563833 403024 563999 403058
rect 564033 403024 564199 403058
rect 564233 403024 564399 403058
rect 564433 403024 564599 403058
rect 564633 403024 564799 403058
rect 564833 403024 564999 403058
rect 565033 403024 565199 403058
rect 565233 403024 565399 403058
rect 565433 403024 565599 403058
rect 565633 403024 565736 403058
rect 560600 402991 565736 403024
rect 560613 358989 560813 359015
rect 560871 358989 561071 359015
rect 561129 358989 561329 359015
rect 561387 358989 561587 359015
rect 561645 358989 561845 359015
rect 561903 358989 562103 359015
rect 562161 358989 562361 359015
rect 562419 358989 562619 359015
rect 562677 358989 562877 359015
rect 562935 358989 563135 359015
rect 563193 358989 563393 359015
rect 563451 358989 563651 359015
rect 563709 358989 563909 359015
rect 563967 358989 564167 359015
rect 564225 358989 564425 359015
rect 564483 358989 564683 359015
rect 564741 358989 564941 359015
rect 564999 358989 565199 359015
rect 565257 358989 565457 359015
rect 565515 358989 565715 359015
rect 574751 358919 574951 358945
rect 575009 358919 575209 358945
rect 575267 358919 575467 358945
rect 575525 358919 575725 358945
rect 575783 358919 575983 358945
rect 576041 358919 576241 358945
rect 576299 358919 576499 358945
rect 576557 358919 576757 358945
rect 576815 358919 577015 358945
rect 577073 358919 577273 358945
rect 577331 358919 577531 358945
rect 577589 358919 577789 358945
rect 577847 358919 578047 358945
rect 578105 358919 578305 358945
rect 578363 358919 578563 358945
rect 578621 358919 578821 358945
rect 578879 358919 579079 358945
rect 579137 358919 579337 358945
rect 579395 358919 579595 358945
rect 579653 358919 579853 358945
rect 560613 357963 560813 357989
rect 560871 357963 561071 357989
rect 561129 357963 561329 357989
rect 561387 357963 561587 357989
rect 561645 357963 561845 357989
rect 561903 357963 562103 357989
rect 562161 357963 562361 357989
rect 562419 357963 562619 357989
rect 562677 357963 562877 357989
rect 562935 357963 563135 357989
rect 563193 357963 563393 357989
rect 563451 357963 563651 357989
rect 563709 357963 563909 357989
rect 563967 357963 564167 357989
rect 564225 357963 564425 357989
rect 564483 357963 564683 357989
rect 564741 357963 564941 357989
rect 564999 357963 565199 357989
rect 565257 357963 565457 357989
rect 565515 357963 565715 357989
rect 560668 357773 560788 357963
rect 560924 357773 561044 357963
rect 561180 357773 561300 357963
rect 561436 357773 561556 357963
rect 561692 357773 561812 357963
rect 561948 357773 562068 357963
rect 562204 357773 562324 357963
rect 562460 357773 562580 357963
rect 562716 357773 562836 357963
rect 562972 357773 563092 357963
rect 563228 357773 563348 357963
rect 563484 357773 563604 357963
rect 563740 357773 563860 357963
rect 563996 357773 564116 357963
rect 564252 357773 564372 357963
rect 564508 357773 564628 357963
rect 564764 357773 564884 357963
rect 565020 357773 565140 357963
rect 565276 357773 565396 357963
rect 565532 357773 565652 357963
rect 574751 357893 574951 357919
rect 575009 357893 575209 357919
rect 575267 357893 575467 357919
rect 575525 357893 575725 357919
rect 575783 357893 575983 357919
rect 576041 357893 576241 357919
rect 576299 357893 576499 357919
rect 576557 357893 576757 357919
rect 576815 357893 577015 357919
rect 577073 357893 577273 357919
rect 577331 357893 577531 357919
rect 577589 357893 577789 357919
rect 577847 357893 578047 357919
rect 578105 357893 578305 357919
rect 578363 357893 578563 357919
rect 578621 357893 578821 357919
rect 578879 357893 579079 357919
rect 579137 357893 579337 357919
rect 579395 357893 579595 357919
rect 579653 357893 579853 357919
rect 560556 357740 565692 357773
rect 560556 357706 560755 357740
rect 560789 357706 560955 357740
rect 560989 357706 561155 357740
rect 561189 357706 561355 357740
rect 561389 357706 561555 357740
rect 561589 357706 561755 357740
rect 561789 357706 561955 357740
rect 561989 357706 562155 357740
rect 562189 357706 562355 357740
rect 562389 357706 562555 357740
rect 562589 357706 562755 357740
rect 562789 357706 562955 357740
rect 562989 357706 563155 357740
rect 563189 357706 563355 357740
rect 563389 357706 563555 357740
rect 563589 357706 563755 357740
rect 563789 357706 563955 357740
rect 563989 357706 564155 357740
rect 564189 357706 564355 357740
rect 564389 357706 564555 357740
rect 564589 357706 564755 357740
rect 564789 357706 564955 357740
rect 564989 357706 565155 357740
rect 565189 357706 565355 357740
rect 565389 357706 565555 357740
rect 565589 357706 565692 357740
rect 560556 357673 565692 357706
rect 574822 357647 574942 357893
rect 575078 357647 575198 357893
rect 575334 357647 575454 357893
rect 575590 357647 575710 357893
rect 575846 357647 575966 357893
rect 576102 357647 576222 357893
rect 576358 357647 576478 357893
rect 576614 357647 576734 357893
rect 576870 357647 576990 357893
rect 577126 357647 577246 357893
rect 577382 357647 577502 357893
rect 577638 357647 577758 357893
rect 577894 357647 578014 357893
rect 578150 357647 578270 357893
rect 578406 357647 578526 357893
rect 578662 357647 578782 357893
rect 578918 357647 579038 357893
rect 579174 357647 579294 357893
rect 579430 357647 579550 357893
rect 579686 357647 579806 357893
rect 574658 357614 579946 357647
rect 574658 357580 574729 357614
rect 574763 357580 574929 357614
rect 574963 357580 575129 357614
rect 575163 357580 575329 357614
rect 575363 357580 575529 357614
rect 575563 357580 575729 357614
rect 575763 357580 575929 357614
rect 575963 357580 576129 357614
rect 576163 357580 576329 357614
rect 576363 357580 576529 357614
rect 576563 357580 576729 357614
rect 576763 357580 576929 357614
rect 576963 357580 577129 357614
rect 577163 357580 577329 357614
rect 577363 357580 577529 357614
rect 577563 357580 577729 357614
rect 577763 357580 577929 357614
rect 577963 357580 578129 357614
rect 578163 357580 578329 357614
rect 578363 357580 578529 357614
rect 578563 357580 578729 357614
rect 578763 357580 578929 357614
rect 578963 357580 579129 357614
rect 579163 357580 579329 357614
rect 579363 357580 579529 357614
rect 579563 357580 579729 357614
rect 579763 357580 579946 357614
rect 574658 357547 579946 357580
rect 575199 312751 575399 312777
rect 575457 312751 575657 312777
rect 575715 312751 575915 312777
rect 575973 312751 576173 312777
rect 576231 312751 576431 312777
rect 576489 312751 576689 312777
rect 576747 312751 576947 312777
rect 577005 312751 577205 312777
rect 577263 312751 577463 312777
rect 577521 312751 577721 312777
rect 577779 312751 577979 312777
rect 578037 312751 578237 312777
rect 578295 312751 578495 312777
rect 578553 312751 578753 312777
rect 578811 312751 579011 312777
rect 579069 312751 579269 312777
rect 579327 312751 579527 312777
rect 579585 312751 579785 312777
rect 579843 312751 580043 312777
rect 580101 312751 580301 312777
rect 560475 312681 560675 312707
rect 560733 312681 560933 312707
rect 560991 312681 561191 312707
rect 561249 312681 561449 312707
rect 561507 312681 561707 312707
rect 561765 312681 561965 312707
rect 562023 312681 562223 312707
rect 562281 312681 562481 312707
rect 562539 312681 562739 312707
rect 562797 312681 562997 312707
rect 563055 312681 563255 312707
rect 563313 312681 563513 312707
rect 563571 312681 563771 312707
rect 563829 312681 564029 312707
rect 564087 312681 564287 312707
rect 564345 312681 564545 312707
rect 564603 312681 564803 312707
rect 564861 312681 565061 312707
rect 565119 312681 565319 312707
rect 565377 312681 565577 312707
rect 575199 311725 575399 311751
rect 575457 311725 575657 311751
rect 575715 311725 575915 311751
rect 575973 311725 576173 311751
rect 576231 311725 576431 311751
rect 576489 311725 576689 311751
rect 576747 311725 576947 311751
rect 577005 311725 577205 311751
rect 577263 311725 577463 311751
rect 577521 311725 577721 311751
rect 577779 311725 577979 311751
rect 578037 311725 578237 311751
rect 578295 311725 578495 311751
rect 578553 311725 578753 311751
rect 578811 311725 579011 311751
rect 579069 311725 579269 311751
rect 579327 311725 579527 311751
rect 579585 311725 579785 311751
rect 579843 311725 580043 311751
rect 580101 311725 580301 311751
rect 560475 311655 560675 311681
rect 560733 311655 560933 311681
rect 560991 311655 561191 311681
rect 561249 311655 561449 311681
rect 561507 311655 561707 311681
rect 561765 311655 561965 311681
rect 562023 311655 562223 311681
rect 562281 311655 562481 311681
rect 562539 311655 562739 311681
rect 562797 311655 562997 311681
rect 563055 311655 563255 311681
rect 563313 311655 563513 311681
rect 563571 311655 563771 311681
rect 563829 311655 564029 311681
rect 564087 311655 564287 311681
rect 564345 311655 564545 311681
rect 564603 311655 564803 311681
rect 564861 311655 565061 311681
rect 565119 311655 565319 311681
rect 565377 311655 565577 311681
rect 560530 311465 560650 311655
rect 560786 311465 560906 311655
rect 561042 311465 561162 311655
rect 561298 311465 561418 311655
rect 561554 311465 561674 311655
rect 561810 311465 561930 311655
rect 562066 311465 562186 311655
rect 562322 311465 562442 311655
rect 562578 311465 562698 311655
rect 562834 311465 562954 311655
rect 563090 311465 563210 311655
rect 563346 311465 563466 311655
rect 563602 311465 563722 311655
rect 563858 311465 563978 311655
rect 564114 311465 564234 311655
rect 564370 311465 564490 311655
rect 564626 311465 564746 311655
rect 564882 311465 565002 311655
rect 565138 311465 565258 311655
rect 565394 311465 565514 311655
rect 575270 311479 575390 311725
rect 575526 311479 575646 311725
rect 575782 311479 575902 311725
rect 576038 311479 576158 311725
rect 576294 311479 576414 311725
rect 576550 311479 576670 311725
rect 576806 311479 576926 311725
rect 577062 311479 577182 311725
rect 577318 311479 577438 311725
rect 577574 311479 577694 311725
rect 577830 311479 577950 311725
rect 578086 311479 578206 311725
rect 578342 311479 578462 311725
rect 578598 311479 578718 311725
rect 578854 311479 578974 311725
rect 579110 311479 579230 311725
rect 579366 311479 579486 311725
rect 579622 311479 579742 311725
rect 579878 311479 579998 311725
rect 580134 311479 580254 311725
rect 560418 311432 565554 311465
rect 560418 311398 560617 311432
rect 560651 311398 560817 311432
rect 560851 311398 561017 311432
rect 561051 311398 561217 311432
rect 561251 311398 561417 311432
rect 561451 311398 561617 311432
rect 561651 311398 561817 311432
rect 561851 311398 562017 311432
rect 562051 311398 562217 311432
rect 562251 311398 562417 311432
rect 562451 311398 562617 311432
rect 562651 311398 562817 311432
rect 562851 311398 563017 311432
rect 563051 311398 563217 311432
rect 563251 311398 563417 311432
rect 563451 311398 563617 311432
rect 563651 311398 563817 311432
rect 563851 311398 564017 311432
rect 564051 311398 564217 311432
rect 564251 311398 564417 311432
rect 564451 311398 564617 311432
rect 564651 311398 564817 311432
rect 564851 311398 565017 311432
rect 565051 311398 565217 311432
rect 565251 311398 565417 311432
rect 565451 311398 565554 311432
rect 560418 311365 565554 311398
rect 575106 311446 580394 311479
rect 575106 311412 575177 311446
rect 575211 311412 575377 311446
rect 575411 311412 575577 311446
rect 575611 311412 575777 311446
rect 575811 311412 575977 311446
rect 576011 311412 576177 311446
rect 576211 311412 576377 311446
rect 576411 311412 576577 311446
rect 576611 311412 576777 311446
rect 576811 311412 576977 311446
rect 577011 311412 577177 311446
rect 577211 311412 577377 311446
rect 577411 311412 577577 311446
rect 577611 311412 577777 311446
rect 577811 311412 577977 311446
rect 578011 311412 578177 311446
rect 578211 311412 578377 311446
rect 578411 311412 578577 311446
rect 578611 311412 578777 311446
rect 578811 311412 578977 311446
rect 579011 311412 579177 311446
rect 579211 311412 579377 311446
rect 579411 311412 579577 311446
rect 579611 311412 579777 311446
rect 579811 311412 579977 311446
rect 580011 311412 580177 311446
rect 580211 311412 580394 311446
rect 575106 311379 580394 311412
<< polycont >>
rect 560863 492166 560897 492200
rect 561063 492166 561097 492200
rect 561263 492166 561297 492200
rect 561463 492166 561497 492200
rect 561663 492166 561697 492200
rect 561863 492166 561897 492200
rect 562063 492166 562097 492200
rect 562263 492166 562297 492200
rect 562463 492166 562497 492200
rect 562663 492166 562697 492200
rect 562863 492166 562897 492200
rect 563063 492166 563097 492200
rect 563263 492166 563297 492200
rect 563463 492166 563497 492200
rect 563663 492166 563697 492200
rect 563863 492166 563897 492200
rect 564063 492166 564097 492200
rect 564263 492166 564297 492200
rect 564463 492166 564497 492200
rect 564663 492166 564697 492200
rect 564863 492166 564897 492200
rect 565063 492166 565097 492200
rect 565263 492166 565297 492200
rect 565463 492166 565497 492200
rect 565663 492166 565697 492200
rect 575255 491884 575289 491918
rect 575455 491884 575489 491918
rect 575655 491884 575689 491918
rect 575855 491884 575889 491918
rect 576055 491884 576089 491918
rect 576255 491884 576289 491918
rect 576455 491884 576489 491918
rect 576655 491884 576689 491918
rect 576855 491884 576889 491918
rect 577055 491884 577089 491918
rect 577255 491884 577289 491918
rect 577455 491884 577489 491918
rect 577655 491884 577689 491918
rect 577855 491884 577889 491918
rect 578055 491884 578089 491918
rect 578255 491884 578289 491918
rect 578455 491884 578489 491918
rect 578655 491884 578689 491918
rect 578855 491884 578889 491918
rect 579055 491884 579089 491918
rect 579255 491884 579289 491918
rect 579455 491884 579489 491918
rect 579655 491884 579689 491918
rect 579855 491884 579889 491918
rect 580055 491884 580089 491918
rect 580255 491884 580289 491918
rect 560799 403024 560833 403058
rect 560999 403024 561033 403058
rect 561199 403024 561233 403058
rect 561399 403024 561433 403058
rect 561599 403024 561633 403058
rect 561799 403024 561833 403058
rect 561999 403024 562033 403058
rect 562199 403024 562233 403058
rect 562399 403024 562433 403058
rect 562599 403024 562633 403058
rect 562799 403024 562833 403058
rect 562999 403024 563033 403058
rect 563199 403024 563233 403058
rect 563399 403024 563433 403058
rect 563599 403024 563633 403058
rect 563799 403024 563833 403058
rect 563999 403024 564033 403058
rect 564199 403024 564233 403058
rect 564399 403024 564433 403058
rect 564599 403024 564633 403058
rect 564799 403024 564833 403058
rect 564999 403024 565033 403058
rect 565199 403024 565233 403058
rect 565399 403024 565433 403058
rect 565599 403024 565633 403058
rect 560755 357706 560789 357740
rect 560955 357706 560989 357740
rect 561155 357706 561189 357740
rect 561355 357706 561389 357740
rect 561555 357706 561589 357740
rect 561755 357706 561789 357740
rect 561955 357706 561989 357740
rect 562155 357706 562189 357740
rect 562355 357706 562389 357740
rect 562555 357706 562589 357740
rect 562755 357706 562789 357740
rect 562955 357706 562989 357740
rect 563155 357706 563189 357740
rect 563355 357706 563389 357740
rect 563555 357706 563589 357740
rect 563755 357706 563789 357740
rect 563955 357706 563989 357740
rect 564155 357706 564189 357740
rect 564355 357706 564389 357740
rect 564555 357706 564589 357740
rect 564755 357706 564789 357740
rect 564955 357706 564989 357740
rect 565155 357706 565189 357740
rect 565355 357706 565389 357740
rect 565555 357706 565589 357740
rect 574729 357580 574763 357614
rect 574929 357580 574963 357614
rect 575129 357580 575163 357614
rect 575329 357580 575363 357614
rect 575529 357580 575563 357614
rect 575729 357580 575763 357614
rect 575929 357580 575963 357614
rect 576129 357580 576163 357614
rect 576329 357580 576363 357614
rect 576529 357580 576563 357614
rect 576729 357580 576763 357614
rect 576929 357580 576963 357614
rect 577129 357580 577163 357614
rect 577329 357580 577363 357614
rect 577529 357580 577563 357614
rect 577729 357580 577763 357614
rect 577929 357580 577963 357614
rect 578129 357580 578163 357614
rect 578329 357580 578363 357614
rect 578529 357580 578563 357614
rect 578729 357580 578763 357614
rect 578929 357580 578963 357614
rect 579129 357580 579163 357614
rect 579329 357580 579363 357614
rect 579529 357580 579563 357614
rect 579729 357580 579763 357614
rect 560617 311398 560651 311432
rect 560817 311398 560851 311432
rect 561017 311398 561051 311432
rect 561217 311398 561251 311432
rect 561417 311398 561451 311432
rect 561617 311398 561651 311432
rect 561817 311398 561851 311432
rect 562017 311398 562051 311432
rect 562217 311398 562251 311432
rect 562417 311398 562451 311432
rect 562617 311398 562651 311432
rect 562817 311398 562851 311432
rect 563017 311398 563051 311432
rect 563217 311398 563251 311432
rect 563417 311398 563451 311432
rect 563617 311398 563651 311432
rect 563817 311398 563851 311432
rect 564017 311398 564051 311432
rect 564217 311398 564251 311432
rect 564417 311398 564451 311432
rect 564617 311398 564651 311432
rect 564817 311398 564851 311432
rect 565017 311398 565051 311432
rect 565217 311398 565251 311432
rect 565417 311398 565451 311432
rect 575177 311412 575211 311446
rect 575377 311412 575411 311446
rect 575577 311412 575611 311446
rect 575777 311412 575811 311446
rect 575977 311412 576011 311446
rect 576177 311412 576211 311446
rect 576377 311412 576411 311446
rect 576577 311412 576611 311446
rect 576777 311412 576811 311446
rect 576977 311412 577011 311446
rect 577177 311412 577211 311446
rect 577377 311412 577411 311446
rect 577577 311412 577611 311446
rect 577777 311412 577811 311446
rect 577977 311412 578011 311446
rect 578177 311412 578211 311446
rect 578377 311412 578411 311446
rect 578577 311412 578611 311446
rect 578777 311412 578811 311446
rect 578977 311412 579011 311446
rect 579177 311412 579211 311446
rect 579377 311412 579411 311446
rect 579577 311412 579611 311446
rect 579777 311412 579811 311446
rect 579977 311412 580011 311446
rect 580177 311412 580211 311446
<< locali >>
rect 560664 493846 565978 493859
rect 560664 493812 560863 493846
rect 560897 493812 561063 493846
rect 561097 493812 561263 493846
rect 561297 493812 561463 493846
rect 561497 493812 561663 493846
rect 561697 493812 561863 493846
rect 561897 493812 562063 493846
rect 562097 493812 562263 493846
rect 562297 493812 562463 493846
rect 562497 493812 562663 493846
rect 562697 493812 562863 493846
rect 562897 493812 563063 493846
rect 563097 493812 563263 493846
rect 563297 493812 563463 493846
rect 563497 493812 563663 493846
rect 563697 493812 563863 493846
rect 563897 493812 564063 493846
rect 564097 493812 564263 493846
rect 564297 493812 564463 493846
rect 564497 493812 564663 493846
rect 564697 493812 564863 493846
rect 564897 493812 565063 493846
rect 565097 493812 565263 493846
rect 565297 493812 565463 493846
rect 565497 493812 565663 493846
rect 565697 493812 565978 493846
rect 560664 493799 565978 493812
rect 560402 493699 560462 493701
rect 560402 493639 565880 493699
rect 560402 492531 560496 493639
rect 560356 492513 560496 492531
rect 560344 492469 560496 492513
rect 560344 492363 560367 492469
rect 560473 492363 560496 492469
rect 560675 493434 560709 493453
rect 560675 493362 560709 493374
rect 560675 493290 560709 493306
rect 560675 493218 560709 493238
rect 560675 493146 560709 493170
rect 560675 493074 560709 493102
rect 560675 493002 560709 493034
rect 560675 492932 560709 492966
rect 560675 492864 560709 492896
rect 560675 492796 560709 492824
rect 560675 492728 560709 492752
rect 560675 492660 560709 492680
rect 560675 492592 560709 492608
rect 560675 492524 560709 492536
rect 560675 492445 560709 492464
rect 560933 493434 560967 493639
rect 560933 493362 560967 493374
rect 560933 493290 560967 493306
rect 560933 493218 560967 493238
rect 560933 493146 560967 493170
rect 560933 493074 560967 493102
rect 560933 493002 560967 493034
rect 560933 492932 560967 492966
rect 560933 492864 560967 492896
rect 560933 492796 560967 492824
rect 560933 492728 560967 492752
rect 560933 492660 560967 492680
rect 560933 492592 560967 492608
rect 560933 492524 560967 492536
rect 560933 492445 560967 492464
rect 561191 493434 561225 493453
rect 561191 493362 561225 493374
rect 561191 493290 561225 493306
rect 561191 493218 561225 493238
rect 561191 493146 561225 493170
rect 561191 493074 561225 493102
rect 561191 493002 561225 493034
rect 561191 492932 561225 492966
rect 561191 492864 561225 492896
rect 561191 492796 561225 492824
rect 561191 492728 561225 492752
rect 561191 492660 561225 492680
rect 561191 492592 561225 492608
rect 561191 492524 561225 492536
rect 561191 492379 561225 492464
rect 561449 493434 561483 493639
rect 561449 493362 561483 493374
rect 561449 493290 561483 493306
rect 561449 493218 561483 493238
rect 561449 493146 561483 493170
rect 561449 493074 561483 493102
rect 561449 493002 561483 493034
rect 561449 492932 561483 492966
rect 561449 492864 561483 492896
rect 561449 492796 561483 492824
rect 561449 492728 561483 492752
rect 561449 492660 561483 492680
rect 561449 492592 561483 492608
rect 561449 492524 561483 492536
rect 561449 492445 561483 492464
rect 561707 493434 561741 493453
rect 561707 493362 561741 493374
rect 561707 493290 561741 493306
rect 561707 493218 561741 493238
rect 561707 493146 561741 493170
rect 561707 493074 561741 493102
rect 561707 493002 561741 493034
rect 561707 492932 561741 492966
rect 561707 492864 561741 492896
rect 561707 492796 561741 492824
rect 561707 492728 561741 492752
rect 561707 492660 561741 492680
rect 561707 492592 561741 492608
rect 561707 492524 561741 492536
rect 561707 492379 561741 492464
rect 561965 493434 561999 493639
rect 561965 493362 561999 493374
rect 561965 493290 561999 493306
rect 561965 493218 561999 493238
rect 561965 493146 561999 493170
rect 561965 493074 561999 493102
rect 561965 493002 561999 493034
rect 561965 492932 561999 492966
rect 561965 492864 561999 492896
rect 561965 492796 561999 492824
rect 561965 492728 561999 492752
rect 561965 492660 561999 492680
rect 561965 492592 561999 492608
rect 561965 492524 561999 492536
rect 561965 492445 561999 492464
rect 562223 493434 562257 493453
rect 562223 493362 562257 493374
rect 562223 493290 562257 493306
rect 562223 493218 562257 493238
rect 562223 493146 562257 493170
rect 562223 493074 562257 493102
rect 562223 493002 562257 493034
rect 562223 492932 562257 492966
rect 562223 492864 562257 492896
rect 562223 492796 562257 492824
rect 562223 492728 562257 492752
rect 562223 492660 562257 492680
rect 562223 492592 562257 492608
rect 562223 492524 562257 492536
rect 562223 492379 562257 492464
rect 562481 493434 562515 493639
rect 562481 493362 562515 493374
rect 562481 493290 562515 493306
rect 562481 493218 562515 493238
rect 562481 493146 562515 493170
rect 562481 493074 562515 493102
rect 562481 493002 562515 493034
rect 562481 492932 562515 492966
rect 562481 492864 562515 492896
rect 562481 492796 562515 492824
rect 562481 492728 562515 492752
rect 562481 492660 562515 492680
rect 562481 492592 562515 492608
rect 562481 492524 562515 492536
rect 562481 492445 562515 492464
rect 562739 493434 562773 493453
rect 562739 493362 562773 493374
rect 562739 493290 562773 493306
rect 562739 493218 562773 493238
rect 562739 493146 562773 493170
rect 562739 493074 562773 493102
rect 562739 493002 562773 493034
rect 562739 492932 562773 492966
rect 562739 492864 562773 492896
rect 562739 492796 562773 492824
rect 562739 492728 562773 492752
rect 562739 492660 562773 492680
rect 562739 492592 562773 492608
rect 562739 492524 562773 492536
rect 562739 492379 562773 492464
rect 562997 493434 563031 493639
rect 562997 493362 563031 493374
rect 562997 493290 563031 493306
rect 562997 493218 563031 493238
rect 562997 493146 563031 493170
rect 562997 493074 563031 493102
rect 562997 493002 563031 493034
rect 562997 492932 563031 492966
rect 562997 492864 563031 492896
rect 562997 492796 563031 492824
rect 562997 492728 563031 492752
rect 562997 492660 563031 492680
rect 562997 492592 563031 492608
rect 562997 492524 563031 492536
rect 562997 492445 563031 492464
rect 563255 493434 563289 493453
rect 563255 493362 563289 493374
rect 563255 493290 563289 493306
rect 563255 493218 563289 493238
rect 563255 493146 563289 493170
rect 563255 493074 563289 493102
rect 563255 493002 563289 493034
rect 563255 492932 563289 492966
rect 563255 492864 563289 492896
rect 563255 492796 563289 492824
rect 563255 492728 563289 492752
rect 563255 492660 563289 492680
rect 563255 492592 563289 492608
rect 563255 492524 563289 492536
rect 563255 492379 563289 492464
rect 563513 493434 563547 493639
rect 563513 493362 563547 493374
rect 563513 493290 563547 493306
rect 563513 493218 563547 493238
rect 563513 493146 563547 493170
rect 563513 493074 563547 493102
rect 563513 493002 563547 493034
rect 563513 492932 563547 492966
rect 563513 492864 563547 492896
rect 563513 492796 563547 492824
rect 563513 492728 563547 492752
rect 563513 492660 563547 492680
rect 563513 492592 563547 492608
rect 563513 492524 563547 492536
rect 563513 492445 563547 492464
rect 563771 493434 563805 493453
rect 563771 493362 563805 493374
rect 563771 493290 563805 493306
rect 563771 493218 563805 493238
rect 563771 493146 563805 493170
rect 563771 493074 563805 493102
rect 563771 493002 563805 493034
rect 563771 492932 563805 492966
rect 563771 492864 563805 492896
rect 563771 492796 563805 492824
rect 563771 492728 563805 492752
rect 563771 492660 563805 492680
rect 563771 492592 563805 492608
rect 563771 492524 563805 492536
rect 563771 492379 563805 492464
rect 564029 493434 564063 493639
rect 564029 493362 564063 493374
rect 564029 493290 564063 493306
rect 564029 493218 564063 493238
rect 564029 493146 564063 493170
rect 564029 493074 564063 493102
rect 564029 493002 564063 493034
rect 564029 492932 564063 492966
rect 564029 492864 564063 492896
rect 564029 492796 564063 492824
rect 564029 492728 564063 492752
rect 564029 492660 564063 492680
rect 564029 492592 564063 492608
rect 564029 492524 564063 492536
rect 564029 492445 564063 492464
rect 564287 493434 564321 493453
rect 564287 493362 564321 493374
rect 564287 493290 564321 493306
rect 564287 493218 564321 493238
rect 564287 493146 564321 493170
rect 564287 493074 564321 493102
rect 564287 493002 564321 493034
rect 564287 492932 564321 492966
rect 564287 492864 564321 492896
rect 564287 492796 564321 492824
rect 564287 492728 564321 492752
rect 564287 492660 564321 492680
rect 564287 492592 564321 492608
rect 564287 492524 564321 492536
rect 564287 492379 564321 492464
rect 564545 493434 564579 493639
rect 564545 493362 564579 493374
rect 564545 493290 564579 493306
rect 564545 493218 564579 493238
rect 564545 493146 564579 493170
rect 564545 493074 564579 493102
rect 564545 493002 564579 493034
rect 564545 492932 564579 492966
rect 564545 492864 564579 492896
rect 564545 492796 564579 492824
rect 564545 492728 564579 492752
rect 564545 492660 564579 492680
rect 564545 492592 564579 492608
rect 564545 492524 564579 492536
rect 564545 492445 564579 492464
rect 564803 493434 564837 493453
rect 564803 493362 564837 493374
rect 564803 493290 564837 493306
rect 564803 493218 564837 493238
rect 564803 493146 564837 493170
rect 564803 493074 564837 493102
rect 564803 493002 564837 493034
rect 564803 492932 564837 492966
rect 564803 492864 564837 492896
rect 564803 492796 564837 492824
rect 564803 492728 564837 492752
rect 564803 492660 564837 492680
rect 564803 492592 564837 492608
rect 564803 492524 564837 492536
rect 564803 492379 564837 492464
rect 565061 493434 565095 493639
rect 565061 493362 565095 493374
rect 565061 493290 565095 493306
rect 565061 493218 565095 493238
rect 565061 493146 565095 493170
rect 565061 493074 565095 493102
rect 565061 493002 565095 493034
rect 565061 492932 565095 492966
rect 565061 492864 565095 492896
rect 565061 492796 565095 492824
rect 565061 492728 565095 492752
rect 565061 492660 565095 492680
rect 565061 492592 565095 492608
rect 565061 492524 565095 492536
rect 565061 492445 565095 492464
rect 565319 493434 565353 493453
rect 565319 493362 565353 493374
rect 565319 493290 565353 493306
rect 565319 493218 565353 493238
rect 565319 493146 565353 493170
rect 565319 493074 565353 493102
rect 565319 493002 565353 493034
rect 565319 492932 565353 492966
rect 565319 492864 565353 492896
rect 565319 492796 565353 492824
rect 565319 492728 565353 492752
rect 565319 492660 565353 492680
rect 565319 492592 565353 492608
rect 565319 492524 565353 492536
rect 565319 492379 565353 492464
rect 565577 493434 565611 493639
rect 575184 493620 580570 493633
rect 575184 493586 575255 493620
rect 575289 493586 575455 493620
rect 575489 493586 575655 493620
rect 575689 493586 575855 493620
rect 575889 493586 576055 493620
rect 576089 493586 576255 493620
rect 576289 493586 576455 493620
rect 576489 493586 576655 493620
rect 576689 493586 576855 493620
rect 576889 493586 577055 493620
rect 577089 493586 577255 493620
rect 577289 493586 577455 493620
rect 577489 493586 577655 493620
rect 577689 493586 577855 493620
rect 577889 493586 578055 493620
rect 578089 493586 578255 493620
rect 578289 493586 578455 493620
rect 578489 493586 578655 493620
rect 578689 493586 578855 493620
rect 578889 493586 579055 493620
rect 579089 493586 579255 493620
rect 579289 493586 579455 493620
rect 579489 493586 579655 493620
rect 579689 493586 579855 493620
rect 579889 493586 580055 493620
rect 580089 493586 580255 493620
rect 580289 493586 580570 493620
rect 575184 493573 580570 493586
rect 576734 493530 576894 493573
rect 576734 493496 576795 493530
rect 576829 493496 576894 493530
rect 576734 493493 576894 493496
rect 578034 493530 578194 493573
rect 578034 493496 578095 493530
rect 578129 493496 578194 493530
rect 578034 493493 578194 493496
rect 579334 493530 579494 493573
rect 579334 493496 579395 493530
rect 579429 493496 579494 493530
rect 579334 493493 579494 493496
rect 580482 493480 580542 493573
rect 574994 493453 575054 493455
rect 565577 493362 565611 493374
rect 565577 493290 565611 493306
rect 565577 493218 565611 493238
rect 565577 493146 565611 493170
rect 565577 493074 565611 493102
rect 565577 493002 565611 493034
rect 565577 492932 565611 492966
rect 565577 492864 565611 492896
rect 565577 492796 565611 492824
rect 565577 492728 565611 492752
rect 565577 492660 565611 492680
rect 565577 492592 565611 492608
rect 565577 492524 565611 492536
rect 565577 492445 565611 492464
rect 565835 493434 565869 493453
rect 565835 493362 565869 493374
rect 565835 493290 565869 493306
rect 565835 493218 565869 493238
rect 565835 493146 565869 493170
rect 565835 493074 565869 493102
rect 565835 493002 565869 493034
rect 565835 492932 565869 492966
rect 565835 492864 565869 492896
rect 565835 492796 565869 492824
rect 565835 492728 565869 492752
rect 565835 492660 565869 492680
rect 565835 492592 565869 492608
rect 565835 492524 565869 492536
rect 565835 492453 565869 492464
rect 574994 493413 580412 493453
rect 580482 493446 580495 493480
rect 580529 493446 580542 493480
rect 574994 493393 580410 493413
rect 565835 492433 565894 492453
rect 566088 492436 566248 492437
rect 566088 492433 566115 492436
rect 565835 492379 566115 492433
rect 560344 492321 560496 492363
rect 560402 492213 560496 492321
rect 560662 492330 566115 492379
rect 566221 492433 566248 492436
rect 566221 492330 566254 492433
rect 560662 492319 566254 492330
rect 560402 492200 565800 492213
rect 560402 492166 560863 492200
rect 560897 492166 561063 492200
rect 561097 492166 561263 492200
rect 561297 492166 561463 492200
rect 561497 492166 561663 492200
rect 561697 492166 561863 492200
rect 561897 492166 562063 492200
rect 562097 492166 562263 492200
rect 562297 492166 562463 492200
rect 562497 492166 562663 492200
rect 562697 492166 562863 492200
rect 562897 492166 563063 492200
rect 563097 492166 563263 492200
rect 563297 492166 563463 492200
rect 563497 492166 563663 492200
rect 563697 492166 563863 492200
rect 563897 492166 564063 492200
rect 564097 492166 564263 492200
rect 564297 492166 564463 492200
rect 564497 492166 564663 492200
rect 564697 492166 564863 492200
rect 564897 492166 565063 492200
rect 565097 492166 565263 492200
rect 565297 492166 565463 492200
rect 565497 492166 565663 492200
rect 565697 492166 565800 492200
rect 560402 492153 565800 492166
rect 565890 492106 565950 492189
rect 562142 492076 562302 492099
rect 562142 492042 562203 492076
rect 562237 492042 562302 492076
rect 562142 491979 562302 492042
rect 563442 492076 563602 492099
rect 563442 492042 563503 492076
rect 563537 492042 563602 492076
rect 563442 491979 563602 492042
rect 564742 492076 564902 492099
rect 564742 492042 564803 492076
rect 564837 492042 564902 492076
rect 564742 491979 564902 492042
rect 565890 492072 565903 492106
rect 565937 492072 565950 492106
rect 565890 491979 565950 492072
rect 574994 492047 575054 493393
rect 575231 493208 575265 493227
rect 575231 493136 575265 493148
rect 575231 493064 575265 493080
rect 575231 492992 575265 493012
rect 575231 492920 575265 492944
rect 575231 492848 575265 492876
rect 575231 492776 575265 492808
rect 575231 492706 575265 492740
rect 575231 492638 575265 492670
rect 575231 492570 575265 492598
rect 575231 492502 575265 492526
rect 575231 492434 575265 492454
rect 575231 492366 575265 492382
rect 575231 492298 575265 492310
rect 575231 492093 575265 492238
rect 575489 493208 575523 493393
rect 575489 493136 575523 493148
rect 575489 493064 575523 493080
rect 575489 492992 575523 493012
rect 575489 492920 575523 492944
rect 575489 492848 575523 492876
rect 575489 492776 575523 492808
rect 575489 492706 575523 492740
rect 575489 492638 575523 492670
rect 575489 492570 575523 492598
rect 575489 492502 575523 492526
rect 575489 492434 575523 492454
rect 575489 492366 575523 492382
rect 575489 492298 575523 492310
rect 575489 492219 575523 492238
rect 575747 493208 575781 493227
rect 575747 493136 575781 493148
rect 575747 493064 575781 493080
rect 575747 492992 575781 493012
rect 575747 492920 575781 492944
rect 575747 492848 575781 492876
rect 575747 492776 575781 492808
rect 575747 492706 575781 492740
rect 575747 492638 575781 492670
rect 575747 492570 575781 492598
rect 575747 492502 575781 492526
rect 575747 492434 575781 492454
rect 575747 492366 575781 492382
rect 575747 492298 575781 492310
rect 575747 492093 575781 492238
rect 576005 493208 576039 493393
rect 576005 493136 576039 493148
rect 576005 493064 576039 493080
rect 576005 492992 576039 493012
rect 576005 492920 576039 492944
rect 576005 492848 576039 492876
rect 576005 492776 576039 492808
rect 576005 492706 576039 492740
rect 576005 492638 576039 492670
rect 576005 492570 576039 492598
rect 576005 492502 576039 492526
rect 576005 492434 576039 492454
rect 576005 492366 576039 492382
rect 576005 492298 576039 492310
rect 576005 492219 576039 492238
rect 576263 493208 576297 493227
rect 576263 493136 576297 493148
rect 576263 493064 576297 493080
rect 576263 492992 576297 493012
rect 576263 492920 576297 492944
rect 576263 492848 576297 492876
rect 576263 492776 576297 492808
rect 576263 492706 576297 492740
rect 576263 492638 576297 492670
rect 576263 492570 576297 492598
rect 576263 492502 576297 492526
rect 576263 492434 576297 492454
rect 576263 492366 576297 492382
rect 576263 492298 576297 492310
rect 576263 492093 576297 492238
rect 576521 493208 576555 493393
rect 576521 493136 576555 493148
rect 576521 493064 576555 493080
rect 576521 492992 576555 493012
rect 576521 492920 576555 492944
rect 576521 492848 576555 492876
rect 576521 492776 576555 492808
rect 576521 492706 576555 492740
rect 576521 492638 576555 492670
rect 576521 492570 576555 492598
rect 576521 492502 576555 492526
rect 576521 492434 576555 492454
rect 576521 492366 576555 492382
rect 576521 492298 576555 492310
rect 576521 492219 576555 492238
rect 576779 493208 576813 493227
rect 576779 493136 576813 493148
rect 576779 493064 576813 493080
rect 576779 492992 576813 493012
rect 576779 492920 576813 492944
rect 576779 492848 576813 492876
rect 576779 492776 576813 492808
rect 576779 492706 576813 492740
rect 576779 492638 576813 492670
rect 576779 492570 576813 492598
rect 576779 492502 576813 492526
rect 576779 492434 576813 492454
rect 576779 492366 576813 492382
rect 576779 492298 576813 492310
rect 576779 492093 576813 492238
rect 577037 493208 577071 493393
rect 577037 493136 577071 493148
rect 577037 493064 577071 493080
rect 577037 492992 577071 493012
rect 577037 492920 577071 492944
rect 577037 492848 577071 492876
rect 577037 492776 577071 492808
rect 577037 492706 577071 492740
rect 577037 492638 577071 492670
rect 577037 492570 577071 492598
rect 577037 492502 577071 492526
rect 577037 492434 577071 492454
rect 577037 492366 577071 492382
rect 577037 492298 577071 492310
rect 577037 492219 577071 492238
rect 577295 493208 577329 493227
rect 577295 493136 577329 493148
rect 577295 493064 577329 493080
rect 577295 492992 577329 493012
rect 577295 492920 577329 492944
rect 577295 492848 577329 492876
rect 577295 492776 577329 492808
rect 577295 492706 577329 492740
rect 577295 492638 577329 492670
rect 577295 492570 577329 492598
rect 577295 492502 577329 492526
rect 577295 492434 577329 492454
rect 577295 492366 577329 492382
rect 577295 492298 577329 492310
rect 577295 492093 577329 492238
rect 577553 493208 577587 493393
rect 577553 493136 577587 493148
rect 577553 493064 577587 493080
rect 577553 492992 577587 493012
rect 577553 492920 577587 492944
rect 577553 492848 577587 492876
rect 577553 492776 577587 492808
rect 577553 492706 577587 492740
rect 577553 492638 577587 492670
rect 577553 492570 577587 492598
rect 577553 492502 577587 492526
rect 577553 492434 577587 492454
rect 577553 492366 577587 492382
rect 577553 492298 577587 492310
rect 577553 492219 577587 492238
rect 577811 493208 577845 493227
rect 577811 493136 577845 493148
rect 577811 493064 577845 493080
rect 577811 492992 577845 493012
rect 577811 492920 577845 492944
rect 577811 492848 577845 492876
rect 577811 492776 577845 492808
rect 577811 492706 577845 492740
rect 577811 492638 577845 492670
rect 577811 492570 577845 492598
rect 577811 492502 577845 492526
rect 577811 492434 577845 492454
rect 577811 492366 577845 492382
rect 577811 492298 577845 492310
rect 577811 492093 577845 492238
rect 578069 493208 578103 493393
rect 578069 493136 578103 493148
rect 578069 493064 578103 493080
rect 578069 492992 578103 493012
rect 578069 492920 578103 492944
rect 578069 492848 578103 492876
rect 578069 492776 578103 492808
rect 578069 492706 578103 492740
rect 578069 492638 578103 492670
rect 578069 492570 578103 492598
rect 578069 492502 578103 492526
rect 578069 492434 578103 492454
rect 578069 492366 578103 492382
rect 578069 492298 578103 492310
rect 578069 492219 578103 492238
rect 578327 493208 578361 493227
rect 578327 493136 578361 493148
rect 578327 493064 578361 493080
rect 578327 492992 578361 493012
rect 578327 492920 578361 492944
rect 578327 492848 578361 492876
rect 578327 492776 578361 492808
rect 578327 492706 578361 492740
rect 578327 492638 578361 492670
rect 578327 492570 578361 492598
rect 578327 492502 578361 492526
rect 578327 492434 578361 492454
rect 578327 492366 578361 492382
rect 578327 492298 578361 492310
rect 578327 492093 578361 492238
rect 578585 493208 578619 493393
rect 578585 493136 578619 493148
rect 578585 493064 578619 493080
rect 578585 492992 578619 493012
rect 578585 492920 578619 492944
rect 578585 492848 578619 492876
rect 578585 492776 578619 492808
rect 578585 492706 578619 492740
rect 578585 492638 578619 492670
rect 578585 492570 578619 492598
rect 578585 492502 578619 492526
rect 578585 492434 578619 492454
rect 578585 492366 578619 492382
rect 578585 492298 578619 492310
rect 578585 492219 578619 492238
rect 578843 493208 578877 493227
rect 578843 493136 578877 493148
rect 578843 493064 578877 493080
rect 578843 492992 578877 493012
rect 578843 492920 578877 492944
rect 578843 492848 578877 492876
rect 578843 492776 578877 492808
rect 578843 492706 578877 492740
rect 578843 492638 578877 492670
rect 578843 492570 578877 492598
rect 578843 492502 578877 492526
rect 578843 492434 578877 492454
rect 578843 492366 578877 492382
rect 578843 492298 578877 492310
rect 578843 492093 578877 492238
rect 579101 493208 579135 493393
rect 579101 493136 579135 493148
rect 579101 493064 579135 493080
rect 579101 492992 579135 493012
rect 579101 492920 579135 492944
rect 579101 492848 579135 492876
rect 579101 492776 579135 492808
rect 579101 492706 579135 492740
rect 579101 492638 579135 492670
rect 579101 492570 579135 492598
rect 579101 492502 579135 492526
rect 579101 492434 579135 492454
rect 579101 492366 579135 492382
rect 579101 492298 579135 492310
rect 579101 492219 579135 492238
rect 579359 493208 579393 493227
rect 579359 493136 579393 493148
rect 579359 493064 579393 493080
rect 579359 492992 579393 493012
rect 579359 492920 579393 492944
rect 579359 492848 579393 492876
rect 579359 492776 579393 492808
rect 579359 492706 579393 492740
rect 579359 492638 579393 492670
rect 579359 492570 579393 492598
rect 579359 492502 579393 492526
rect 579359 492434 579393 492454
rect 579359 492366 579393 492382
rect 579359 492298 579393 492310
rect 579359 492093 579393 492238
rect 579617 493208 579651 493393
rect 579617 493136 579651 493148
rect 579617 493064 579651 493080
rect 579617 492992 579651 493012
rect 579617 492920 579651 492944
rect 579617 492848 579651 492876
rect 579617 492776 579651 492808
rect 579617 492706 579651 492740
rect 579617 492638 579651 492670
rect 579617 492570 579651 492598
rect 579617 492502 579651 492526
rect 579617 492434 579651 492454
rect 579617 492366 579651 492382
rect 579617 492298 579651 492310
rect 579617 492219 579651 492238
rect 579875 493208 579909 493227
rect 579875 493136 579909 493148
rect 579875 493064 579909 493080
rect 579875 492992 579909 493012
rect 579875 492920 579909 492944
rect 579875 492848 579909 492876
rect 579875 492776 579909 492808
rect 579875 492706 579909 492740
rect 579875 492638 579909 492670
rect 579875 492570 579909 492598
rect 579875 492502 579909 492526
rect 579875 492434 579909 492454
rect 579875 492366 579909 492382
rect 579875 492298 579909 492310
rect 579875 492093 579909 492238
rect 580133 493208 580167 493393
rect 580482 493363 580542 493446
rect 580133 493136 580167 493148
rect 580133 493064 580167 493080
rect 580133 492992 580167 493012
rect 580133 492920 580167 492944
rect 580133 492848 580167 492876
rect 580133 492776 580167 492808
rect 580133 492706 580167 492740
rect 580133 492638 580167 492670
rect 580133 492570 580167 492598
rect 580133 492502 580167 492526
rect 580133 492434 580167 492454
rect 580133 492366 580167 492382
rect 580133 492298 580167 492310
rect 580133 492219 580167 492238
rect 580391 493208 580425 493227
rect 580391 493136 580425 493148
rect 580391 493064 580425 493080
rect 580391 492992 580425 493012
rect 580391 492920 580425 492944
rect 580391 492848 580425 492876
rect 580391 492776 580425 492808
rect 580391 492706 580425 492740
rect 580391 492638 580425 492670
rect 580391 492570 580425 492598
rect 580391 492502 580425 492526
rect 580391 492434 580425 492454
rect 580391 492366 580425 492382
rect 580391 492298 580425 492310
rect 580391 492217 580425 492238
rect 580428 492100 580656 492137
rect 580428 492093 580584 492100
rect 560664 491966 565978 491979
rect 560664 491932 560863 491966
rect 560897 491932 561063 491966
rect 561097 491932 561263 491966
rect 561297 491932 561463 491966
rect 561497 491932 561663 491966
rect 561697 491932 561863 491966
rect 561897 491932 562063 491966
rect 562097 491932 562263 491966
rect 562297 491932 562463 491966
rect 562497 491932 562663 491966
rect 562697 491932 562863 491966
rect 562897 491932 563063 491966
rect 563097 491932 563263 491966
rect 563297 491932 563463 491966
rect 563497 491932 563663 491966
rect 563697 491932 563863 491966
rect 563897 491932 564063 491966
rect 564097 491932 564263 491966
rect 564297 491932 564463 491966
rect 564497 491932 564663 491966
rect 564697 491932 564863 491966
rect 564897 491932 565063 491966
rect 565097 491932 565263 491966
rect 565297 491932 565463 491966
rect 565497 491932 565663 491966
rect 565697 491932 565978 491966
rect 560664 491919 565978 491932
rect 574938 491958 575054 492047
rect 575178 492066 580584 492093
rect 580618 492066 580656 492100
rect 575178 492033 580656 492066
rect 574938 491924 574977 491958
rect 575011 491931 575054 491958
rect 575011 491924 580472 491931
rect 574938 491918 580472 491924
rect 574938 491884 575255 491918
rect 575289 491884 575455 491918
rect 575489 491884 575655 491918
rect 575689 491884 575855 491918
rect 575889 491884 576055 491918
rect 576089 491884 576255 491918
rect 576289 491884 576455 491918
rect 576489 491884 576655 491918
rect 576689 491884 576855 491918
rect 576889 491884 577055 491918
rect 577089 491884 577255 491918
rect 577289 491884 577455 491918
rect 577489 491884 577655 491918
rect 577689 491884 577855 491918
rect 577889 491884 578055 491918
rect 578089 491884 578255 491918
rect 578289 491884 578455 491918
rect 578489 491884 578655 491918
rect 578689 491884 578855 491918
rect 578889 491884 579055 491918
rect 579089 491884 579255 491918
rect 579289 491884 579455 491918
rect 579489 491884 579655 491918
rect 579689 491884 579855 491918
rect 579889 491884 580055 491918
rect 580089 491884 580255 491918
rect 580289 491884 580472 491918
rect 574938 491873 580472 491884
rect 574976 491871 580472 491873
rect 575184 491740 580570 491753
rect 575184 491706 575255 491740
rect 575289 491706 575455 491740
rect 575489 491706 575655 491740
rect 575689 491706 575855 491740
rect 575889 491706 576055 491740
rect 576089 491706 576255 491740
rect 576289 491706 576455 491740
rect 576489 491706 576655 491740
rect 576689 491706 576855 491740
rect 576889 491706 577055 491740
rect 577089 491706 577255 491740
rect 577289 491706 577455 491740
rect 577489 491706 577655 491740
rect 577689 491706 577855 491740
rect 577889 491706 578055 491740
rect 578089 491706 578255 491740
rect 578289 491706 578455 491740
rect 578489 491706 578655 491740
rect 578689 491706 578855 491740
rect 578889 491706 579055 491740
rect 579089 491706 579255 491740
rect 579289 491706 579455 491740
rect 579489 491706 579655 491740
rect 579689 491706 579855 491740
rect 579889 491706 580055 491740
rect 580089 491706 580255 491740
rect 580289 491706 580570 491740
rect 575184 491693 580570 491706
rect 560600 404704 565914 404717
rect 560600 404670 560799 404704
rect 560833 404670 560999 404704
rect 561033 404670 561199 404704
rect 561233 404670 561399 404704
rect 561433 404670 561599 404704
rect 561633 404670 561799 404704
rect 561833 404670 561999 404704
rect 562033 404670 562199 404704
rect 562233 404670 562399 404704
rect 562433 404670 562599 404704
rect 562633 404670 562799 404704
rect 562833 404670 562999 404704
rect 563033 404670 563199 404704
rect 563233 404670 563399 404704
rect 563433 404670 563599 404704
rect 563633 404670 563799 404704
rect 563833 404670 563999 404704
rect 564033 404670 564199 404704
rect 564233 404670 564399 404704
rect 564433 404670 564599 404704
rect 564633 404670 564799 404704
rect 564833 404670 564999 404704
rect 565033 404670 565199 404704
rect 565233 404670 565399 404704
rect 565433 404670 565599 404704
rect 565633 404670 565914 404704
rect 560600 404657 565914 404670
rect 560338 404557 560398 404559
rect 560338 404497 565816 404557
rect 560338 403389 560432 404497
rect 560292 403371 560432 403389
rect 560280 403327 560432 403371
rect 560280 403221 560303 403327
rect 560409 403221 560432 403327
rect 560611 404292 560645 404311
rect 560611 404220 560645 404232
rect 560611 404148 560645 404164
rect 560611 404076 560645 404096
rect 560611 404004 560645 404028
rect 560611 403932 560645 403960
rect 560611 403860 560645 403892
rect 560611 403790 560645 403824
rect 560611 403722 560645 403754
rect 560611 403654 560645 403682
rect 560611 403586 560645 403610
rect 560611 403518 560645 403538
rect 560611 403450 560645 403466
rect 560611 403382 560645 403394
rect 560611 403303 560645 403322
rect 560869 404292 560903 404497
rect 560869 404220 560903 404232
rect 560869 404148 560903 404164
rect 560869 404076 560903 404096
rect 560869 404004 560903 404028
rect 560869 403932 560903 403960
rect 560869 403860 560903 403892
rect 560869 403790 560903 403824
rect 560869 403722 560903 403754
rect 560869 403654 560903 403682
rect 560869 403586 560903 403610
rect 560869 403518 560903 403538
rect 560869 403450 560903 403466
rect 560869 403382 560903 403394
rect 560869 403303 560903 403322
rect 561127 404292 561161 404311
rect 561127 404220 561161 404232
rect 561127 404148 561161 404164
rect 561127 404076 561161 404096
rect 561127 404004 561161 404028
rect 561127 403932 561161 403960
rect 561127 403860 561161 403892
rect 561127 403790 561161 403824
rect 561127 403722 561161 403754
rect 561127 403654 561161 403682
rect 561127 403586 561161 403610
rect 561127 403518 561161 403538
rect 561127 403450 561161 403466
rect 561127 403382 561161 403394
rect 561127 403237 561161 403322
rect 561385 404292 561419 404497
rect 561385 404220 561419 404232
rect 561385 404148 561419 404164
rect 561385 404076 561419 404096
rect 561385 404004 561419 404028
rect 561385 403932 561419 403960
rect 561385 403860 561419 403892
rect 561385 403790 561419 403824
rect 561385 403722 561419 403754
rect 561385 403654 561419 403682
rect 561385 403586 561419 403610
rect 561385 403518 561419 403538
rect 561385 403450 561419 403466
rect 561385 403382 561419 403394
rect 561385 403303 561419 403322
rect 561643 404292 561677 404311
rect 561643 404220 561677 404232
rect 561643 404148 561677 404164
rect 561643 404076 561677 404096
rect 561643 404004 561677 404028
rect 561643 403932 561677 403960
rect 561643 403860 561677 403892
rect 561643 403790 561677 403824
rect 561643 403722 561677 403754
rect 561643 403654 561677 403682
rect 561643 403586 561677 403610
rect 561643 403518 561677 403538
rect 561643 403450 561677 403466
rect 561643 403382 561677 403394
rect 561643 403237 561677 403322
rect 561901 404292 561935 404497
rect 561901 404220 561935 404232
rect 561901 404148 561935 404164
rect 561901 404076 561935 404096
rect 561901 404004 561935 404028
rect 561901 403932 561935 403960
rect 561901 403860 561935 403892
rect 561901 403790 561935 403824
rect 561901 403722 561935 403754
rect 561901 403654 561935 403682
rect 561901 403586 561935 403610
rect 561901 403518 561935 403538
rect 561901 403450 561935 403466
rect 561901 403382 561935 403394
rect 561901 403303 561935 403322
rect 562159 404292 562193 404311
rect 562159 404220 562193 404232
rect 562159 404148 562193 404164
rect 562159 404076 562193 404096
rect 562159 404004 562193 404028
rect 562159 403932 562193 403960
rect 562159 403860 562193 403892
rect 562159 403790 562193 403824
rect 562159 403722 562193 403754
rect 562159 403654 562193 403682
rect 562159 403586 562193 403610
rect 562159 403518 562193 403538
rect 562159 403450 562193 403466
rect 562159 403382 562193 403394
rect 562159 403237 562193 403322
rect 562417 404292 562451 404497
rect 562417 404220 562451 404232
rect 562417 404148 562451 404164
rect 562417 404076 562451 404096
rect 562417 404004 562451 404028
rect 562417 403932 562451 403960
rect 562417 403860 562451 403892
rect 562417 403790 562451 403824
rect 562417 403722 562451 403754
rect 562417 403654 562451 403682
rect 562417 403586 562451 403610
rect 562417 403518 562451 403538
rect 562417 403450 562451 403466
rect 562417 403382 562451 403394
rect 562417 403303 562451 403322
rect 562675 404292 562709 404311
rect 562675 404220 562709 404232
rect 562675 404148 562709 404164
rect 562675 404076 562709 404096
rect 562675 404004 562709 404028
rect 562675 403932 562709 403960
rect 562675 403860 562709 403892
rect 562675 403790 562709 403824
rect 562675 403722 562709 403754
rect 562675 403654 562709 403682
rect 562675 403586 562709 403610
rect 562675 403518 562709 403538
rect 562675 403450 562709 403466
rect 562675 403382 562709 403394
rect 562675 403237 562709 403322
rect 562933 404292 562967 404497
rect 562933 404220 562967 404232
rect 562933 404148 562967 404164
rect 562933 404076 562967 404096
rect 562933 404004 562967 404028
rect 562933 403932 562967 403960
rect 562933 403860 562967 403892
rect 562933 403790 562967 403824
rect 562933 403722 562967 403754
rect 562933 403654 562967 403682
rect 562933 403586 562967 403610
rect 562933 403518 562967 403538
rect 562933 403450 562967 403466
rect 562933 403382 562967 403394
rect 562933 403303 562967 403322
rect 563191 404292 563225 404311
rect 563191 404220 563225 404232
rect 563191 404148 563225 404164
rect 563191 404076 563225 404096
rect 563191 404004 563225 404028
rect 563191 403932 563225 403960
rect 563191 403860 563225 403892
rect 563191 403790 563225 403824
rect 563191 403722 563225 403754
rect 563191 403654 563225 403682
rect 563191 403586 563225 403610
rect 563191 403518 563225 403538
rect 563191 403450 563225 403466
rect 563191 403382 563225 403394
rect 563191 403237 563225 403322
rect 563449 404292 563483 404497
rect 563449 404220 563483 404232
rect 563449 404148 563483 404164
rect 563449 404076 563483 404096
rect 563449 404004 563483 404028
rect 563449 403932 563483 403960
rect 563449 403860 563483 403892
rect 563449 403790 563483 403824
rect 563449 403722 563483 403754
rect 563449 403654 563483 403682
rect 563449 403586 563483 403610
rect 563449 403518 563483 403538
rect 563449 403450 563483 403466
rect 563449 403382 563483 403394
rect 563449 403303 563483 403322
rect 563707 404292 563741 404311
rect 563707 404220 563741 404232
rect 563707 404148 563741 404164
rect 563707 404076 563741 404096
rect 563707 404004 563741 404028
rect 563707 403932 563741 403960
rect 563707 403860 563741 403892
rect 563707 403790 563741 403824
rect 563707 403722 563741 403754
rect 563707 403654 563741 403682
rect 563707 403586 563741 403610
rect 563707 403518 563741 403538
rect 563707 403450 563741 403466
rect 563707 403382 563741 403394
rect 563707 403237 563741 403322
rect 563965 404292 563999 404497
rect 563965 404220 563999 404232
rect 563965 404148 563999 404164
rect 563965 404076 563999 404096
rect 563965 404004 563999 404028
rect 563965 403932 563999 403960
rect 563965 403860 563999 403892
rect 563965 403790 563999 403824
rect 563965 403722 563999 403754
rect 563965 403654 563999 403682
rect 563965 403586 563999 403610
rect 563965 403518 563999 403538
rect 563965 403450 563999 403466
rect 563965 403382 563999 403394
rect 563965 403303 563999 403322
rect 564223 404292 564257 404311
rect 564223 404220 564257 404232
rect 564223 404148 564257 404164
rect 564223 404076 564257 404096
rect 564223 404004 564257 404028
rect 564223 403932 564257 403960
rect 564223 403860 564257 403892
rect 564223 403790 564257 403824
rect 564223 403722 564257 403754
rect 564223 403654 564257 403682
rect 564223 403586 564257 403610
rect 564223 403518 564257 403538
rect 564223 403450 564257 403466
rect 564223 403382 564257 403394
rect 564223 403237 564257 403322
rect 564481 404292 564515 404497
rect 564481 404220 564515 404232
rect 564481 404148 564515 404164
rect 564481 404076 564515 404096
rect 564481 404004 564515 404028
rect 564481 403932 564515 403960
rect 564481 403860 564515 403892
rect 564481 403790 564515 403824
rect 564481 403722 564515 403754
rect 564481 403654 564515 403682
rect 564481 403586 564515 403610
rect 564481 403518 564515 403538
rect 564481 403450 564515 403466
rect 564481 403382 564515 403394
rect 564481 403303 564515 403322
rect 564739 404292 564773 404311
rect 564739 404220 564773 404232
rect 564739 404148 564773 404164
rect 564739 404076 564773 404096
rect 564739 404004 564773 404028
rect 564739 403932 564773 403960
rect 564739 403860 564773 403892
rect 564739 403790 564773 403824
rect 564739 403722 564773 403754
rect 564739 403654 564773 403682
rect 564739 403586 564773 403610
rect 564739 403518 564773 403538
rect 564739 403450 564773 403466
rect 564739 403382 564773 403394
rect 564739 403237 564773 403322
rect 564997 404292 565031 404497
rect 564997 404220 565031 404232
rect 564997 404148 565031 404164
rect 564997 404076 565031 404096
rect 564997 404004 565031 404028
rect 564997 403932 565031 403960
rect 564997 403860 565031 403892
rect 564997 403790 565031 403824
rect 564997 403722 565031 403754
rect 564997 403654 565031 403682
rect 564997 403586 565031 403610
rect 564997 403518 565031 403538
rect 564997 403450 565031 403466
rect 564997 403382 565031 403394
rect 564997 403303 565031 403322
rect 565255 404292 565289 404311
rect 565255 404220 565289 404232
rect 565255 404148 565289 404164
rect 565255 404076 565289 404096
rect 565255 404004 565289 404028
rect 565255 403932 565289 403960
rect 565255 403860 565289 403892
rect 565255 403790 565289 403824
rect 565255 403722 565289 403754
rect 565255 403654 565289 403682
rect 565255 403586 565289 403610
rect 565255 403518 565289 403538
rect 565255 403450 565289 403466
rect 565255 403382 565289 403394
rect 565255 403237 565289 403322
rect 565513 404292 565547 404497
rect 565513 404220 565547 404232
rect 565513 404148 565547 404164
rect 565513 404076 565547 404096
rect 565513 404004 565547 404028
rect 565513 403932 565547 403960
rect 565513 403860 565547 403892
rect 565513 403790 565547 403824
rect 565513 403722 565547 403754
rect 565513 403654 565547 403682
rect 565513 403586 565547 403610
rect 565513 403518 565547 403538
rect 565513 403450 565547 403466
rect 565513 403382 565547 403394
rect 565513 403303 565547 403322
rect 565771 404292 565805 404311
rect 565771 404220 565805 404232
rect 565771 404148 565805 404164
rect 565771 404076 565805 404096
rect 565771 404004 565805 404028
rect 565771 403932 565805 403960
rect 565771 403860 565805 403892
rect 565771 403790 565805 403824
rect 565771 403722 565805 403754
rect 565771 403654 565805 403682
rect 565771 403586 565805 403610
rect 565771 403518 565805 403538
rect 565771 403450 565805 403466
rect 565771 403382 565805 403394
rect 565771 403311 565805 403322
rect 565771 403291 565830 403311
rect 566024 403294 566184 403295
rect 566024 403291 566051 403294
rect 565771 403237 566051 403291
rect 560280 403179 560432 403221
rect 560338 403071 560432 403179
rect 560598 403188 566051 403237
rect 566157 403291 566184 403294
rect 566157 403188 566190 403291
rect 560598 403177 566190 403188
rect 560338 403058 565736 403071
rect 560338 403024 560799 403058
rect 560833 403024 560999 403058
rect 561033 403024 561199 403058
rect 561233 403024 561399 403058
rect 561433 403024 561599 403058
rect 561633 403024 561799 403058
rect 561833 403024 561999 403058
rect 562033 403024 562199 403058
rect 562233 403024 562399 403058
rect 562433 403024 562599 403058
rect 562633 403024 562799 403058
rect 562833 403024 562999 403058
rect 563033 403024 563199 403058
rect 563233 403024 563399 403058
rect 563433 403024 563599 403058
rect 563633 403024 563799 403058
rect 563833 403024 563999 403058
rect 564033 403024 564199 403058
rect 564233 403024 564399 403058
rect 564433 403024 564599 403058
rect 564633 403024 564799 403058
rect 564833 403024 564999 403058
rect 565033 403024 565199 403058
rect 565233 403024 565399 403058
rect 565433 403024 565599 403058
rect 565633 403024 565736 403058
rect 560338 403011 565736 403024
rect 565826 402964 565886 403047
rect 562078 402934 562238 402957
rect 562078 402900 562139 402934
rect 562173 402900 562238 402934
rect 562078 402837 562238 402900
rect 563378 402934 563538 402957
rect 563378 402900 563439 402934
rect 563473 402900 563538 402934
rect 563378 402837 563538 402900
rect 564678 402934 564838 402957
rect 564678 402900 564739 402934
rect 564773 402900 564838 402934
rect 564678 402837 564838 402900
rect 565826 402930 565839 402964
rect 565873 402930 565886 402964
rect 565826 402837 565886 402930
rect 560600 402824 565914 402837
rect 560600 402790 560799 402824
rect 560833 402790 560999 402824
rect 561033 402790 561199 402824
rect 561233 402790 561399 402824
rect 561433 402790 561599 402824
rect 561633 402790 561799 402824
rect 561833 402790 561999 402824
rect 562033 402790 562199 402824
rect 562233 402790 562399 402824
rect 562433 402790 562599 402824
rect 562633 402790 562799 402824
rect 562833 402790 562999 402824
rect 563033 402790 563199 402824
rect 563233 402790 563399 402824
rect 563433 402790 563599 402824
rect 563633 402790 563799 402824
rect 563833 402790 563999 402824
rect 564033 402790 564199 402824
rect 564233 402790 564399 402824
rect 564433 402790 564599 402824
rect 564633 402790 564799 402824
rect 564833 402790 564999 402824
rect 565033 402790 565199 402824
rect 565233 402790 565399 402824
rect 565433 402790 565599 402824
rect 565633 402790 565914 402824
rect 560600 402777 565914 402790
rect 560556 359386 565870 359399
rect 560556 359352 560755 359386
rect 560789 359352 560955 359386
rect 560989 359352 561155 359386
rect 561189 359352 561355 359386
rect 561389 359352 561555 359386
rect 561589 359352 561755 359386
rect 561789 359352 561955 359386
rect 561989 359352 562155 359386
rect 562189 359352 562355 359386
rect 562389 359352 562555 359386
rect 562589 359352 562755 359386
rect 562789 359352 562955 359386
rect 562989 359352 563155 359386
rect 563189 359352 563355 359386
rect 563389 359352 563555 359386
rect 563589 359352 563755 359386
rect 563789 359352 563955 359386
rect 563989 359352 564155 359386
rect 564189 359352 564355 359386
rect 564389 359352 564555 359386
rect 564589 359352 564755 359386
rect 564789 359352 564955 359386
rect 564989 359352 565155 359386
rect 565189 359352 565355 359386
rect 565389 359352 565555 359386
rect 565589 359352 565870 359386
rect 560556 359339 565870 359352
rect 574658 359316 580044 359329
rect 574658 359282 574729 359316
rect 574763 359282 574929 359316
rect 574963 359282 575129 359316
rect 575163 359282 575329 359316
rect 575363 359282 575529 359316
rect 575563 359282 575729 359316
rect 575763 359282 575929 359316
rect 575963 359282 576129 359316
rect 576163 359282 576329 359316
rect 576363 359282 576529 359316
rect 576563 359282 576729 359316
rect 576763 359282 576929 359316
rect 576963 359282 577129 359316
rect 577163 359282 577329 359316
rect 577363 359282 577529 359316
rect 577563 359282 577729 359316
rect 577763 359282 577929 359316
rect 577963 359282 578129 359316
rect 578163 359282 578329 359316
rect 578363 359282 578529 359316
rect 578563 359282 578729 359316
rect 578763 359282 578929 359316
rect 578963 359282 579129 359316
rect 579163 359282 579329 359316
rect 579363 359282 579529 359316
rect 579563 359282 579729 359316
rect 579763 359282 580044 359316
rect 574658 359269 580044 359282
rect 560294 359239 560354 359241
rect 560294 359179 565772 359239
rect 576208 359226 576368 359269
rect 576208 359192 576269 359226
rect 576303 359192 576368 359226
rect 576208 359189 576368 359192
rect 577508 359226 577668 359269
rect 577508 359192 577569 359226
rect 577603 359192 577668 359226
rect 577508 359189 577668 359192
rect 578808 359226 578968 359269
rect 578808 359192 578869 359226
rect 578903 359192 578968 359226
rect 578808 359189 578968 359192
rect 560294 358071 560388 359179
rect 560248 358053 560388 358071
rect 560236 358009 560388 358053
rect 560236 357903 560259 358009
rect 560365 357903 560388 358009
rect 560567 358974 560601 358993
rect 560567 358902 560601 358914
rect 560567 358830 560601 358846
rect 560567 358758 560601 358778
rect 560567 358686 560601 358710
rect 560567 358614 560601 358642
rect 560567 358542 560601 358574
rect 560567 358472 560601 358506
rect 560567 358404 560601 358436
rect 560567 358336 560601 358364
rect 560567 358268 560601 358292
rect 560567 358200 560601 358220
rect 560567 358132 560601 358148
rect 560567 358064 560601 358076
rect 560567 357985 560601 358004
rect 560825 358974 560859 359179
rect 560825 358902 560859 358914
rect 560825 358830 560859 358846
rect 560825 358758 560859 358778
rect 560825 358686 560859 358710
rect 560825 358614 560859 358642
rect 560825 358542 560859 358574
rect 560825 358472 560859 358506
rect 560825 358404 560859 358436
rect 560825 358336 560859 358364
rect 560825 358268 560859 358292
rect 560825 358200 560859 358220
rect 560825 358132 560859 358148
rect 560825 358064 560859 358076
rect 560825 357985 560859 358004
rect 561083 358974 561117 358993
rect 561083 358902 561117 358914
rect 561083 358830 561117 358846
rect 561083 358758 561117 358778
rect 561083 358686 561117 358710
rect 561083 358614 561117 358642
rect 561083 358542 561117 358574
rect 561083 358472 561117 358506
rect 561083 358404 561117 358436
rect 561083 358336 561117 358364
rect 561083 358268 561117 358292
rect 561083 358200 561117 358220
rect 561083 358132 561117 358148
rect 561083 358064 561117 358076
rect 561083 357919 561117 358004
rect 561341 358974 561375 359179
rect 561341 358902 561375 358914
rect 561341 358830 561375 358846
rect 561341 358758 561375 358778
rect 561341 358686 561375 358710
rect 561341 358614 561375 358642
rect 561341 358542 561375 358574
rect 561341 358472 561375 358506
rect 561341 358404 561375 358436
rect 561341 358336 561375 358364
rect 561341 358268 561375 358292
rect 561341 358200 561375 358220
rect 561341 358132 561375 358148
rect 561341 358064 561375 358076
rect 561341 357985 561375 358004
rect 561599 358974 561633 358993
rect 561599 358902 561633 358914
rect 561599 358830 561633 358846
rect 561599 358758 561633 358778
rect 561599 358686 561633 358710
rect 561599 358614 561633 358642
rect 561599 358542 561633 358574
rect 561599 358472 561633 358506
rect 561599 358404 561633 358436
rect 561599 358336 561633 358364
rect 561599 358268 561633 358292
rect 561599 358200 561633 358220
rect 561599 358132 561633 358148
rect 561599 358064 561633 358076
rect 561599 357919 561633 358004
rect 561857 358974 561891 359179
rect 561857 358902 561891 358914
rect 561857 358830 561891 358846
rect 561857 358758 561891 358778
rect 561857 358686 561891 358710
rect 561857 358614 561891 358642
rect 561857 358542 561891 358574
rect 561857 358472 561891 358506
rect 561857 358404 561891 358436
rect 561857 358336 561891 358364
rect 561857 358268 561891 358292
rect 561857 358200 561891 358220
rect 561857 358132 561891 358148
rect 561857 358064 561891 358076
rect 561857 357985 561891 358004
rect 562115 358974 562149 358993
rect 562115 358902 562149 358914
rect 562115 358830 562149 358846
rect 562115 358758 562149 358778
rect 562115 358686 562149 358710
rect 562115 358614 562149 358642
rect 562115 358542 562149 358574
rect 562115 358472 562149 358506
rect 562115 358404 562149 358436
rect 562115 358336 562149 358364
rect 562115 358268 562149 358292
rect 562115 358200 562149 358220
rect 562115 358132 562149 358148
rect 562115 358064 562149 358076
rect 562115 357919 562149 358004
rect 562373 358974 562407 359179
rect 562373 358902 562407 358914
rect 562373 358830 562407 358846
rect 562373 358758 562407 358778
rect 562373 358686 562407 358710
rect 562373 358614 562407 358642
rect 562373 358542 562407 358574
rect 562373 358472 562407 358506
rect 562373 358404 562407 358436
rect 562373 358336 562407 358364
rect 562373 358268 562407 358292
rect 562373 358200 562407 358220
rect 562373 358132 562407 358148
rect 562373 358064 562407 358076
rect 562373 357985 562407 358004
rect 562631 358974 562665 358993
rect 562631 358902 562665 358914
rect 562631 358830 562665 358846
rect 562631 358758 562665 358778
rect 562631 358686 562665 358710
rect 562631 358614 562665 358642
rect 562631 358542 562665 358574
rect 562631 358472 562665 358506
rect 562631 358404 562665 358436
rect 562631 358336 562665 358364
rect 562631 358268 562665 358292
rect 562631 358200 562665 358220
rect 562631 358132 562665 358148
rect 562631 358064 562665 358076
rect 562631 357919 562665 358004
rect 562889 358974 562923 359179
rect 562889 358902 562923 358914
rect 562889 358830 562923 358846
rect 562889 358758 562923 358778
rect 562889 358686 562923 358710
rect 562889 358614 562923 358642
rect 562889 358542 562923 358574
rect 562889 358472 562923 358506
rect 562889 358404 562923 358436
rect 562889 358336 562923 358364
rect 562889 358268 562923 358292
rect 562889 358200 562923 358220
rect 562889 358132 562923 358148
rect 562889 358064 562923 358076
rect 562889 357985 562923 358004
rect 563147 358974 563181 358993
rect 563147 358902 563181 358914
rect 563147 358830 563181 358846
rect 563147 358758 563181 358778
rect 563147 358686 563181 358710
rect 563147 358614 563181 358642
rect 563147 358542 563181 358574
rect 563147 358472 563181 358506
rect 563147 358404 563181 358436
rect 563147 358336 563181 358364
rect 563147 358268 563181 358292
rect 563147 358200 563181 358220
rect 563147 358132 563181 358148
rect 563147 358064 563181 358076
rect 563147 357919 563181 358004
rect 563405 358974 563439 359179
rect 563405 358902 563439 358914
rect 563405 358830 563439 358846
rect 563405 358758 563439 358778
rect 563405 358686 563439 358710
rect 563405 358614 563439 358642
rect 563405 358542 563439 358574
rect 563405 358472 563439 358506
rect 563405 358404 563439 358436
rect 563405 358336 563439 358364
rect 563405 358268 563439 358292
rect 563405 358200 563439 358220
rect 563405 358132 563439 358148
rect 563405 358064 563439 358076
rect 563405 357985 563439 358004
rect 563663 358974 563697 358993
rect 563663 358902 563697 358914
rect 563663 358830 563697 358846
rect 563663 358758 563697 358778
rect 563663 358686 563697 358710
rect 563663 358614 563697 358642
rect 563663 358542 563697 358574
rect 563663 358472 563697 358506
rect 563663 358404 563697 358436
rect 563663 358336 563697 358364
rect 563663 358268 563697 358292
rect 563663 358200 563697 358220
rect 563663 358132 563697 358148
rect 563663 358064 563697 358076
rect 563663 357919 563697 358004
rect 563921 358974 563955 359179
rect 563921 358902 563955 358914
rect 563921 358830 563955 358846
rect 563921 358758 563955 358778
rect 563921 358686 563955 358710
rect 563921 358614 563955 358642
rect 563921 358542 563955 358574
rect 563921 358472 563955 358506
rect 563921 358404 563955 358436
rect 563921 358336 563955 358364
rect 563921 358268 563955 358292
rect 563921 358200 563955 358220
rect 563921 358132 563955 358148
rect 563921 358064 563955 358076
rect 563921 357985 563955 358004
rect 564179 358974 564213 358993
rect 564179 358902 564213 358914
rect 564179 358830 564213 358846
rect 564179 358758 564213 358778
rect 564179 358686 564213 358710
rect 564179 358614 564213 358642
rect 564179 358542 564213 358574
rect 564179 358472 564213 358506
rect 564179 358404 564213 358436
rect 564179 358336 564213 358364
rect 564179 358268 564213 358292
rect 564179 358200 564213 358220
rect 564179 358132 564213 358148
rect 564179 358064 564213 358076
rect 564179 357919 564213 358004
rect 564437 358974 564471 359179
rect 564437 358902 564471 358914
rect 564437 358830 564471 358846
rect 564437 358758 564471 358778
rect 564437 358686 564471 358710
rect 564437 358614 564471 358642
rect 564437 358542 564471 358574
rect 564437 358472 564471 358506
rect 564437 358404 564471 358436
rect 564437 358336 564471 358364
rect 564437 358268 564471 358292
rect 564437 358200 564471 358220
rect 564437 358132 564471 358148
rect 564437 358064 564471 358076
rect 564437 357985 564471 358004
rect 564695 358974 564729 358993
rect 564695 358902 564729 358914
rect 564695 358830 564729 358846
rect 564695 358758 564729 358778
rect 564695 358686 564729 358710
rect 564695 358614 564729 358642
rect 564695 358542 564729 358574
rect 564695 358472 564729 358506
rect 564695 358404 564729 358436
rect 564695 358336 564729 358364
rect 564695 358268 564729 358292
rect 564695 358200 564729 358220
rect 564695 358132 564729 358148
rect 564695 358064 564729 358076
rect 564695 357919 564729 358004
rect 564953 358974 564987 359179
rect 564953 358902 564987 358914
rect 564953 358830 564987 358846
rect 564953 358758 564987 358778
rect 564953 358686 564987 358710
rect 564953 358614 564987 358642
rect 564953 358542 564987 358574
rect 564953 358472 564987 358506
rect 564953 358404 564987 358436
rect 564953 358336 564987 358364
rect 564953 358268 564987 358292
rect 564953 358200 564987 358220
rect 564953 358132 564987 358148
rect 564953 358064 564987 358076
rect 564953 357985 564987 358004
rect 565211 358974 565245 358993
rect 565211 358902 565245 358914
rect 565211 358830 565245 358846
rect 565211 358758 565245 358778
rect 565211 358686 565245 358710
rect 565211 358614 565245 358642
rect 565211 358542 565245 358574
rect 565211 358472 565245 358506
rect 565211 358404 565245 358436
rect 565211 358336 565245 358364
rect 565211 358268 565245 358292
rect 565211 358200 565245 358220
rect 565211 358132 565245 358148
rect 565211 358064 565245 358076
rect 565211 357919 565245 358004
rect 565469 358974 565503 359179
rect 579956 359176 580016 359269
rect 574468 359149 574528 359151
rect 574468 359109 579886 359149
rect 579956 359142 579969 359176
rect 580003 359142 580016 359176
rect 574468 359089 579884 359109
rect 565469 358902 565503 358914
rect 565469 358830 565503 358846
rect 565469 358758 565503 358778
rect 565469 358686 565503 358710
rect 565469 358614 565503 358642
rect 565469 358542 565503 358574
rect 565469 358472 565503 358506
rect 565469 358404 565503 358436
rect 565469 358336 565503 358364
rect 565469 358268 565503 358292
rect 565469 358200 565503 358220
rect 565469 358132 565503 358148
rect 565469 358064 565503 358076
rect 565469 357985 565503 358004
rect 565727 358974 565761 358993
rect 565727 358902 565761 358914
rect 565727 358830 565761 358846
rect 565727 358758 565761 358778
rect 565727 358686 565761 358710
rect 565727 358614 565761 358642
rect 565727 358542 565761 358574
rect 565727 358472 565761 358506
rect 565727 358404 565761 358436
rect 565727 358336 565761 358364
rect 565727 358268 565761 358292
rect 565727 358200 565761 358220
rect 565727 358132 565761 358148
rect 565727 358064 565761 358076
rect 565727 357993 565761 358004
rect 565727 357973 565786 357993
rect 565980 357976 566140 357977
rect 565980 357973 566007 357976
rect 565727 357919 566007 357973
rect 560236 357861 560388 357903
rect 560294 357753 560388 357861
rect 560554 357870 566007 357919
rect 566113 357973 566140 357976
rect 566113 357870 566146 357973
rect 560554 357859 566146 357870
rect 560294 357740 565692 357753
rect 574468 357743 574528 359089
rect 574705 358904 574739 358923
rect 574705 358832 574739 358844
rect 574705 358760 574739 358776
rect 574705 358688 574739 358708
rect 574705 358616 574739 358640
rect 574705 358544 574739 358572
rect 574705 358472 574739 358504
rect 574705 358402 574739 358436
rect 574705 358334 574739 358366
rect 574705 358266 574739 358294
rect 574705 358198 574739 358222
rect 574705 358130 574739 358150
rect 574705 358062 574739 358078
rect 574705 357994 574739 358006
rect 574705 357789 574739 357934
rect 574963 358904 574997 359089
rect 574963 358832 574997 358844
rect 574963 358760 574997 358776
rect 574963 358688 574997 358708
rect 574963 358616 574997 358640
rect 574963 358544 574997 358572
rect 574963 358472 574997 358504
rect 574963 358402 574997 358436
rect 574963 358334 574997 358366
rect 574963 358266 574997 358294
rect 574963 358198 574997 358222
rect 574963 358130 574997 358150
rect 574963 358062 574997 358078
rect 574963 357994 574997 358006
rect 574963 357915 574997 357934
rect 575221 358904 575255 358923
rect 575221 358832 575255 358844
rect 575221 358760 575255 358776
rect 575221 358688 575255 358708
rect 575221 358616 575255 358640
rect 575221 358544 575255 358572
rect 575221 358472 575255 358504
rect 575221 358402 575255 358436
rect 575221 358334 575255 358366
rect 575221 358266 575255 358294
rect 575221 358198 575255 358222
rect 575221 358130 575255 358150
rect 575221 358062 575255 358078
rect 575221 357994 575255 358006
rect 575221 357789 575255 357934
rect 575479 358904 575513 359089
rect 575479 358832 575513 358844
rect 575479 358760 575513 358776
rect 575479 358688 575513 358708
rect 575479 358616 575513 358640
rect 575479 358544 575513 358572
rect 575479 358472 575513 358504
rect 575479 358402 575513 358436
rect 575479 358334 575513 358366
rect 575479 358266 575513 358294
rect 575479 358198 575513 358222
rect 575479 358130 575513 358150
rect 575479 358062 575513 358078
rect 575479 357994 575513 358006
rect 575479 357915 575513 357934
rect 575737 358904 575771 358923
rect 575737 358832 575771 358844
rect 575737 358760 575771 358776
rect 575737 358688 575771 358708
rect 575737 358616 575771 358640
rect 575737 358544 575771 358572
rect 575737 358472 575771 358504
rect 575737 358402 575771 358436
rect 575737 358334 575771 358366
rect 575737 358266 575771 358294
rect 575737 358198 575771 358222
rect 575737 358130 575771 358150
rect 575737 358062 575771 358078
rect 575737 357994 575771 358006
rect 575737 357789 575771 357934
rect 575995 358904 576029 359089
rect 575995 358832 576029 358844
rect 575995 358760 576029 358776
rect 575995 358688 576029 358708
rect 575995 358616 576029 358640
rect 575995 358544 576029 358572
rect 575995 358472 576029 358504
rect 575995 358402 576029 358436
rect 575995 358334 576029 358366
rect 575995 358266 576029 358294
rect 575995 358198 576029 358222
rect 575995 358130 576029 358150
rect 575995 358062 576029 358078
rect 575995 357994 576029 358006
rect 575995 357915 576029 357934
rect 576253 358904 576287 358923
rect 576253 358832 576287 358844
rect 576253 358760 576287 358776
rect 576253 358688 576287 358708
rect 576253 358616 576287 358640
rect 576253 358544 576287 358572
rect 576253 358472 576287 358504
rect 576253 358402 576287 358436
rect 576253 358334 576287 358366
rect 576253 358266 576287 358294
rect 576253 358198 576287 358222
rect 576253 358130 576287 358150
rect 576253 358062 576287 358078
rect 576253 357994 576287 358006
rect 576253 357789 576287 357934
rect 576511 358904 576545 359089
rect 576511 358832 576545 358844
rect 576511 358760 576545 358776
rect 576511 358688 576545 358708
rect 576511 358616 576545 358640
rect 576511 358544 576545 358572
rect 576511 358472 576545 358504
rect 576511 358402 576545 358436
rect 576511 358334 576545 358366
rect 576511 358266 576545 358294
rect 576511 358198 576545 358222
rect 576511 358130 576545 358150
rect 576511 358062 576545 358078
rect 576511 357994 576545 358006
rect 576511 357915 576545 357934
rect 576769 358904 576803 358923
rect 576769 358832 576803 358844
rect 576769 358760 576803 358776
rect 576769 358688 576803 358708
rect 576769 358616 576803 358640
rect 576769 358544 576803 358572
rect 576769 358472 576803 358504
rect 576769 358402 576803 358436
rect 576769 358334 576803 358366
rect 576769 358266 576803 358294
rect 576769 358198 576803 358222
rect 576769 358130 576803 358150
rect 576769 358062 576803 358078
rect 576769 357994 576803 358006
rect 576769 357789 576803 357934
rect 577027 358904 577061 359089
rect 577027 358832 577061 358844
rect 577027 358760 577061 358776
rect 577027 358688 577061 358708
rect 577027 358616 577061 358640
rect 577027 358544 577061 358572
rect 577027 358472 577061 358504
rect 577027 358402 577061 358436
rect 577027 358334 577061 358366
rect 577027 358266 577061 358294
rect 577027 358198 577061 358222
rect 577027 358130 577061 358150
rect 577027 358062 577061 358078
rect 577027 357994 577061 358006
rect 577027 357915 577061 357934
rect 577285 358904 577319 358923
rect 577285 358832 577319 358844
rect 577285 358760 577319 358776
rect 577285 358688 577319 358708
rect 577285 358616 577319 358640
rect 577285 358544 577319 358572
rect 577285 358472 577319 358504
rect 577285 358402 577319 358436
rect 577285 358334 577319 358366
rect 577285 358266 577319 358294
rect 577285 358198 577319 358222
rect 577285 358130 577319 358150
rect 577285 358062 577319 358078
rect 577285 357994 577319 358006
rect 577285 357789 577319 357934
rect 577543 358904 577577 359089
rect 577543 358832 577577 358844
rect 577543 358760 577577 358776
rect 577543 358688 577577 358708
rect 577543 358616 577577 358640
rect 577543 358544 577577 358572
rect 577543 358472 577577 358504
rect 577543 358402 577577 358436
rect 577543 358334 577577 358366
rect 577543 358266 577577 358294
rect 577543 358198 577577 358222
rect 577543 358130 577577 358150
rect 577543 358062 577577 358078
rect 577543 357994 577577 358006
rect 577543 357915 577577 357934
rect 577801 358904 577835 358923
rect 577801 358832 577835 358844
rect 577801 358760 577835 358776
rect 577801 358688 577835 358708
rect 577801 358616 577835 358640
rect 577801 358544 577835 358572
rect 577801 358472 577835 358504
rect 577801 358402 577835 358436
rect 577801 358334 577835 358366
rect 577801 358266 577835 358294
rect 577801 358198 577835 358222
rect 577801 358130 577835 358150
rect 577801 358062 577835 358078
rect 577801 357994 577835 358006
rect 577801 357789 577835 357934
rect 578059 358904 578093 359089
rect 578059 358832 578093 358844
rect 578059 358760 578093 358776
rect 578059 358688 578093 358708
rect 578059 358616 578093 358640
rect 578059 358544 578093 358572
rect 578059 358472 578093 358504
rect 578059 358402 578093 358436
rect 578059 358334 578093 358366
rect 578059 358266 578093 358294
rect 578059 358198 578093 358222
rect 578059 358130 578093 358150
rect 578059 358062 578093 358078
rect 578059 357994 578093 358006
rect 578059 357915 578093 357934
rect 578317 358904 578351 358923
rect 578317 358832 578351 358844
rect 578317 358760 578351 358776
rect 578317 358688 578351 358708
rect 578317 358616 578351 358640
rect 578317 358544 578351 358572
rect 578317 358472 578351 358504
rect 578317 358402 578351 358436
rect 578317 358334 578351 358366
rect 578317 358266 578351 358294
rect 578317 358198 578351 358222
rect 578317 358130 578351 358150
rect 578317 358062 578351 358078
rect 578317 357994 578351 358006
rect 578317 357789 578351 357934
rect 578575 358904 578609 359089
rect 578575 358832 578609 358844
rect 578575 358760 578609 358776
rect 578575 358688 578609 358708
rect 578575 358616 578609 358640
rect 578575 358544 578609 358572
rect 578575 358472 578609 358504
rect 578575 358402 578609 358436
rect 578575 358334 578609 358366
rect 578575 358266 578609 358294
rect 578575 358198 578609 358222
rect 578575 358130 578609 358150
rect 578575 358062 578609 358078
rect 578575 357994 578609 358006
rect 578575 357915 578609 357934
rect 578833 358904 578867 358923
rect 578833 358832 578867 358844
rect 578833 358760 578867 358776
rect 578833 358688 578867 358708
rect 578833 358616 578867 358640
rect 578833 358544 578867 358572
rect 578833 358472 578867 358504
rect 578833 358402 578867 358436
rect 578833 358334 578867 358366
rect 578833 358266 578867 358294
rect 578833 358198 578867 358222
rect 578833 358130 578867 358150
rect 578833 358062 578867 358078
rect 578833 357994 578867 358006
rect 578833 357789 578867 357934
rect 579091 358904 579125 359089
rect 579091 358832 579125 358844
rect 579091 358760 579125 358776
rect 579091 358688 579125 358708
rect 579091 358616 579125 358640
rect 579091 358544 579125 358572
rect 579091 358472 579125 358504
rect 579091 358402 579125 358436
rect 579091 358334 579125 358366
rect 579091 358266 579125 358294
rect 579091 358198 579125 358222
rect 579091 358130 579125 358150
rect 579091 358062 579125 358078
rect 579091 357994 579125 358006
rect 579091 357915 579125 357934
rect 579349 358904 579383 358923
rect 579349 358832 579383 358844
rect 579349 358760 579383 358776
rect 579349 358688 579383 358708
rect 579349 358616 579383 358640
rect 579349 358544 579383 358572
rect 579349 358472 579383 358504
rect 579349 358402 579383 358436
rect 579349 358334 579383 358366
rect 579349 358266 579383 358294
rect 579349 358198 579383 358222
rect 579349 358130 579383 358150
rect 579349 358062 579383 358078
rect 579349 357994 579383 358006
rect 579349 357789 579383 357934
rect 579607 358904 579641 359089
rect 579956 359059 580016 359142
rect 579607 358832 579641 358844
rect 579607 358760 579641 358776
rect 579607 358688 579641 358708
rect 579607 358616 579641 358640
rect 579607 358544 579641 358572
rect 579607 358472 579641 358504
rect 579607 358402 579641 358436
rect 579607 358334 579641 358366
rect 579607 358266 579641 358294
rect 579607 358198 579641 358222
rect 579607 358130 579641 358150
rect 579607 358062 579641 358078
rect 579607 357994 579641 358006
rect 579607 357915 579641 357934
rect 579865 358904 579899 358923
rect 579865 358832 579899 358844
rect 579865 358760 579899 358776
rect 579865 358688 579899 358708
rect 579865 358616 579899 358640
rect 579865 358544 579899 358572
rect 579865 358472 579899 358504
rect 579865 358402 579899 358436
rect 579865 358334 579899 358366
rect 579865 358266 579899 358294
rect 579865 358198 579899 358222
rect 579865 358130 579899 358150
rect 579865 358062 579899 358078
rect 579865 357994 579899 358006
rect 579865 357913 579899 357934
rect 579902 357796 580130 357833
rect 579902 357789 580058 357796
rect 560294 357706 560755 357740
rect 560789 357706 560955 357740
rect 560989 357706 561155 357740
rect 561189 357706 561355 357740
rect 561389 357706 561555 357740
rect 561589 357706 561755 357740
rect 561789 357706 561955 357740
rect 561989 357706 562155 357740
rect 562189 357706 562355 357740
rect 562389 357706 562555 357740
rect 562589 357706 562755 357740
rect 562789 357706 562955 357740
rect 562989 357706 563155 357740
rect 563189 357706 563355 357740
rect 563389 357706 563555 357740
rect 563589 357706 563755 357740
rect 563789 357706 563955 357740
rect 563989 357706 564155 357740
rect 564189 357706 564355 357740
rect 564389 357706 564555 357740
rect 564589 357706 564755 357740
rect 564789 357706 564955 357740
rect 564989 357706 565155 357740
rect 565189 357706 565355 357740
rect 565389 357706 565555 357740
rect 565589 357706 565692 357740
rect 560294 357693 565692 357706
rect 565782 357646 565842 357729
rect 562034 357616 562194 357639
rect 562034 357582 562095 357616
rect 562129 357582 562194 357616
rect 562034 357519 562194 357582
rect 563334 357616 563494 357639
rect 563334 357582 563395 357616
rect 563429 357582 563494 357616
rect 563334 357519 563494 357582
rect 564634 357616 564794 357639
rect 564634 357582 564695 357616
rect 564729 357582 564794 357616
rect 564634 357519 564794 357582
rect 565782 357612 565795 357646
rect 565829 357612 565842 357646
rect 565782 357519 565842 357612
rect 574412 357654 574528 357743
rect 574652 357762 580058 357789
rect 580092 357762 580130 357796
rect 574652 357729 580130 357762
rect 574412 357620 574451 357654
rect 574485 357627 574528 357654
rect 574485 357620 579946 357627
rect 574412 357614 579946 357620
rect 574412 357580 574729 357614
rect 574763 357580 574929 357614
rect 574963 357580 575129 357614
rect 575163 357580 575329 357614
rect 575363 357580 575529 357614
rect 575563 357580 575729 357614
rect 575763 357580 575929 357614
rect 575963 357580 576129 357614
rect 576163 357580 576329 357614
rect 576363 357580 576529 357614
rect 576563 357580 576729 357614
rect 576763 357580 576929 357614
rect 576963 357580 577129 357614
rect 577163 357580 577329 357614
rect 577363 357580 577529 357614
rect 577563 357580 577729 357614
rect 577763 357580 577929 357614
rect 577963 357580 578129 357614
rect 578163 357580 578329 357614
rect 578363 357580 578529 357614
rect 578563 357580 578729 357614
rect 578763 357580 578929 357614
rect 578963 357580 579129 357614
rect 579163 357580 579329 357614
rect 579363 357580 579529 357614
rect 579563 357580 579729 357614
rect 579763 357580 579946 357614
rect 574412 357569 579946 357580
rect 574450 357567 579946 357569
rect 560556 357506 565870 357519
rect 560556 357472 560755 357506
rect 560789 357472 560955 357506
rect 560989 357472 561155 357506
rect 561189 357472 561355 357506
rect 561389 357472 561555 357506
rect 561589 357472 561755 357506
rect 561789 357472 561955 357506
rect 561989 357472 562155 357506
rect 562189 357472 562355 357506
rect 562389 357472 562555 357506
rect 562589 357472 562755 357506
rect 562789 357472 562955 357506
rect 562989 357472 563155 357506
rect 563189 357472 563355 357506
rect 563389 357472 563555 357506
rect 563589 357472 563755 357506
rect 563789 357472 563955 357506
rect 563989 357472 564155 357506
rect 564189 357472 564355 357506
rect 564389 357472 564555 357506
rect 564589 357472 564755 357506
rect 564789 357472 564955 357506
rect 564989 357472 565155 357506
rect 565189 357472 565355 357506
rect 565389 357472 565555 357506
rect 565589 357472 565870 357506
rect 560556 357459 565870 357472
rect 574658 357436 580044 357449
rect 574658 357402 574729 357436
rect 574763 357402 574929 357436
rect 574963 357402 575129 357436
rect 575163 357402 575329 357436
rect 575363 357402 575529 357436
rect 575563 357402 575729 357436
rect 575763 357402 575929 357436
rect 575963 357402 576129 357436
rect 576163 357402 576329 357436
rect 576363 357402 576529 357436
rect 576563 357402 576729 357436
rect 576763 357402 576929 357436
rect 576963 357402 577129 357436
rect 577163 357402 577329 357436
rect 577363 357402 577529 357436
rect 577563 357402 577729 357436
rect 577763 357402 577929 357436
rect 577963 357402 578129 357436
rect 578163 357402 578329 357436
rect 578363 357402 578529 357436
rect 578563 357402 578729 357436
rect 578763 357402 578929 357436
rect 578963 357402 579129 357436
rect 579163 357402 579329 357436
rect 579363 357402 579529 357436
rect 579563 357402 579729 357436
rect 579763 357402 580044 357436
rect 574658 357389 580044 357402
rect 575106 313148 580492 313161
rect 575106 313114 575177 313148
rect 575211 313114 575377 313148
rect 575411 313114 575577 313148
rect 575611 313114 575777 313148
rect 575811 313114 575977 313148
rect 576011 313114 576177 313148
rect 576211 313114 576377 313148
rect 576411 313114 576577 313148
rect 576611 313114 576777 313148
rect 576811 313114 576977 313148
rect 577011 313114 577177 313148
rect 577211 313114 577377 313148
rect 577411 313114 577577 313148
rect 577611 313114 577777 313148
rect 577811 313114 577977 313148
rect 578011 313114 578177 313148
rect 578211 313114 578377 313148
rect 578411 313114 578577 313148
rect 578611 313114 578777 313148
rect 578811 313114 578977 313148
rect 579011 313114 579177 313148
rect 579211 313114 579377 313148
rect 579411 313114 579577 313148
rect 579611 313114 579777 313148
rect 579811 313114 579977 313148
rect 580011 313114 580177 313148
rect 580211 313114 580492 313148
rect 575106 313101 580492 313114
rect 560418 313078 565732 313091
rect 560418 313044 560617 313078
rect 560651 313044 560817 313078
rect 560851 313044 561017 313078
rect 561051 313044 561217 313078
rect 561251 313044 561417 313078
rect 561451 313044 561617 313078
rect 561651 313044 561817 313078
rect 561851 313044 562017 313078
rect 562051 313044 562217 313078
rect 562251 313044 562417 313078
rect 562451 313044 562617 313078
rect 562651 313044 562817 313078
rect 562851 313044 563017 313078
rect 563051 313044 563217 313078
rect 563251 313044 563417 313078
rect 563451 313044 563617 313078
rect 563651 313044 563817 313078
rect 563851 313044 564017 313078
rect 564051 313044 564217 313078
rect 564251 313044 564417 313078
rect 564451 313044 564617 313078
rect 564651 313044 564817 313078
rect 564851 313044 565017 313078
rect 565051 313044 565217 313078
rect 565251 313044 565417 313078
rect 565451 313044 565732 313078
rect 560418 313031 565732 313044
rect 576656 313058 576816 313101
rect 576656 313024 576717 313058
rect 576751 313024 576816 313058
rect 576656 313021 576816 313024
rect 577956 313058 578116 313101
rect 577956 313024 578017 313058
rect 578051 313024 578116 313058
rect 577956 313021 578116 313024
rect 579256 313058 579416 313101
rect 579256 313024 579317 313058
rect 579351 313024 579416 313058
rect 579256 313021 579416 313024
rect 580404 313008 580464 313101
rect 574916 312981 574976 312983
rect 574916 312941 580334 312981
rect 580404 312974 580417 313008
rect 580451 312974 580464 313008
rect 560156 312931 560216 312933
rect 560156 312871 565634 312931
rect 574916 312921 580332 312941
rect 560156 311763 560250 312871
rect 560110 311745 560250 311763
rect 560098 311701 560250 311745
rect 560098 311595 560121 311701
rect 560227 311595 560250 311701
rect 560429 312666 560463 312685
rect 560429 312594 560463 312606
rect 560429 312522 560463 312538
rect 560429 312450 560463 312470
rect 560429 312378 560463 312402
rect 560429 312306 560463 312334
rect 560429 312234 560463 312266
rect 560429 312164 560463 312198
rect 560429 312096 560463 312128
rect 560429 312028 560463 312056
rect 560429 311960 560463 311984
rect 560429 311892 560463 311912
rect 560429 311824 560463 311840
rect 560429 311756 560463 311768
rect 560429 311677 560463 311696
rect 560687 312666 560721 312871
rect 560687 312594 560721 312606
rect 560687 312522 560721 312538
rect 560687 312450 560721 312470
rect 560687 312378 560721 312402
rect 560687 312306 560721 312334
rect 560687 312234 560721 312266
rect 560687 312164 560721 312198
rect 560687 312096 560721 312128
rect 560687 312028 560721 312056
rect 560687 311960 560721 311984
rect 560687 311892 560721 311912
rect 560687 311824 560721 311840
rect 560687 311756 560721 311768
rect 560687 311677 560721 311696
rect 560945 312666 560979 312685
rect 560945 312594 560979 312606
rect 560945 312522 560979 312538
rect 560945 312450 560979 312470
rect 560945 312378 560979 312402
rect 560945 312306 560979 312334
rect 560945 312234 560979 312266
rect 560945 312164 560979 312198
rect 560945 312096 560979 312128
rect 560945 312028 560979 312056
rect 560945 311960 560979 311984
rect 560945 311892 560979 311912
rect 560945 311824 560979 311840
rect 560945 311756 560979 311768
rect 560945 311611 560979 311696
rect 561203 312666 561237 312871
rect 561203 312594 561237 312606
rect 561203 312522 561237 312538
rect 561203 312450 561237 312470
rect 561203 312378 561237 312402
rect 561203 312306 561237 312334
rect 561203 312234 561237 312266
rect 561203 312164 561237 312198
rect 561203 312096 561237 312128
rect 561203 312028 561237 312056
rect 561203 311960 561237 311984
rect 561203 311892 561237 311912
rect 561203 311824 561237 311840
rect 561203 311756 561237 311768
rect 561203 311677 561237 311696
rect 561461 312666 561495 312685
rect 561461 312594 561495 312606
rect 561461 312522 561495 312538
rect 561461 312450 561495 312470
rect 561461 312378 561495 312402
rect 561461 312306 561495 312334
rect 561461 312234 561495 312266
rect 561461 312164 561495 312198
rect 561461 312096 561495 312128
rect 561461 312028 561495 312056
rect 561461 311960 561495 311984
rect 561461 311892 561495 311912
rect 561461 311824 561495 311840
rect 561461 311756 561495 311768
rect 561461 311611 561495 311696
rect 561719 312666 561753 312871
rect 561719 312594 561753 312606
rect 561719 312522 561753 312538
rect 561719 312450 561753 312470
rect 561719 312378 561753 312402
rect 561719 312306 561753 312334
rect 561719 312234 561753 312266
rect 561719 312164 561753 312198
rect 561719 312096 561753 312128
rect 561719 312028 561753 312056
rect 561719 311960 561753 311984
rect 561719 311892 561753 311912
rect 561719 311824 561753 311840
rect 561719 311756 561753 311768
rect 561719 311677 561753 311696
rect 561977 312666 562011 312685
rect 561977 312594 562011 312606
rect 561977 312522 562011 312538
rect 561977 312450 562011 312470
rect 561977 312378 562011 312402
rect 561977 312306 562011 312334
rect 561977 312234 562011 312266
rect 561977 312164 562011 312198
rect 561977 312096 562011 312128
rect 561977 312028 562011 312056
rect 561977 311960 562011 311984
rect 561977 311892 562011 311912
rect 561977 311824 562011 311840
rect 561977 311756 562011 311768
rect 561977 311611 562011 311696
rect 562235 312666 562269 312871
rect 562235 312594 562269 312606
rect 562235 312522 562269 312538
rect 562235 312450 562269 312470
rect 562235 312378 562269 312402
rect 562235 312306 562269 312334
rect 562235 312234 562269 312266
rect 562235 312164 562269 312198
rect 562235 312096 562269 312128
rect 562235 312028 562269 312056
rect 562235 311960 562269 311984
rect 562235 311892 562269 311912
rect 562235 311824 562269 311840
rect 562235 311756 562269 311768
rect 562235 311677 562269 311696
rect 562493 312666 562527 312685
rect 562493 312594 562527 312606
rect 562493 312522 562527 312538
rect 562493 312450 562527 312470
rect 562493 312378 562527 312402
rect 562493 312306 562527 312334
rect 562493 312234 562527 312266
rect 562493 312164 562527 312198
rect 562493 312096 562527 312128
rect 562493 312028 562527 312056
rect 562493 311960 562527 311984
rect 562493 311892 562527 311912
rect 562493 311824 562527 311840
rect 562493 311756 562527 311768
rect 562493 311611 562527 311696
rect 562751 312666 562785 312871
rect 562751 312594 562785 312606
rect 562751 312522 562785 312538
rect 562751 312450 562785 312470
rect 562751 312378 562785 312402
rect 562751 312306 562785 312334
rect 562751 312234 562785 312266
rect 562751 312164 562785 312198
rect 562751 312096 562785 312128
rect 562751 312028 562785 312056
rect 562751 311960 562785 311984
rect 562751 311892 562785 311912
rect 562751 311824 562785 311840
rect 562751 311756 562785 311768
rect 562751 311677 562785 311696
rect 563009 312666 563043 312685
rect 563009 312594 563043 312606
rect 563009 312522 563043 312538
rect 563009 312450 563043 312470
rect 563009 312378 563043 312402
rect 563009 312306 563043 312334
rect 563009 312234 563043 312266
rect 563009 312164 563043 312198
rect 563009 312096 563043 312128
rect 563009 312028 563043 312056
rect 563009 311960 563043 311984
rect 563009 311892 563043 311912
rect 563009 311824 563043 311840
rect 563009 311756 563043 311768
rect 563009 311611 563043 311696
rect 563267 312666 563301 312871
rect 563267 312594 563301 312606
rect 563267 312522 563301 312538
rect 563267 312450 563301 312470
rect 563267 312378 563301 312402
rect 563267 312306 563301 312334
rect 563267 312234 563301 312266
rect 563267 312164 563301 312198
rect 563267 312096 563301 312128
rect 563267 312028 563301 312056
rect 563267 311960 563301 311984
rect 563267 311892 563301 311912
rect 563267 311824 563301 311840
rect 563267 311756 563301 311768
rect 563267 311677 563301 311696
rect 563525 312666 563559 312685
rect 563525 312594 563559 312606
rect 563525 312522 563559 312538
rect 563525 312450 563559 312470
rect 563525 312378 563559 312402
rect 563525 312306 563559 312334
rect 563525 312234 563559 312266
rect 563525 312164 563559 312198
rect 563525 312096 563559 312128
rect 563525 312028 563559 312056
rect 563525 311960 563559 311984
rect 563525 311892 563559 311912
rect 563525 311824 563559 311840
rect 563525 311756 563559 311768
rect 563525 311611 563559 311696
rect 563783 312666 563817 312871
rect 563783 312594 563817 312606
rect 563783 312522 563817 312538
rect 563783 312450 563817 312470
rect 563783 312378 563817 312402
rect 563783 312306 563817 312334
rect 563783 312234 563817 312266
rect 563783 312164 563817 312198
rect 563783 312096 563817 312128
rect 563783 312028 563817 312056
rect 563783 311960 563817 311984
rect 563783 311892 563817 311912
rect 563783 311824 563817 311840
rect 563783 311756 563817 311768
rect 563783 311677 563817 311696
rect 564041 312666 564075 312685
rect 564041 312594 564075 312606
rect 564041 312522 564075 312538
rect 564041 312450 564075 312470
rect 564041 312378 564075 312402
rect 564041 312306 564075 312334
rect 564041 312234 564075 312266
rect 564041 312164 564075 312198
rect 564041 312096 564075 312128
rect 564041 312028 564075 312056
rect 564041 311960 564075 311984
rect 564041 311892 564075 311912
rect 564041 311824 564075 311840
rect 564041 311756 564075 311768
rect 564041 311611 564075 311696
rect 564299 312666 564333 312871
rect 564299 312594 564333 312606
rect 564299 312522 564333 312538
rect 564299 312450 564333 312470
rect 564299 312378 564333 312402
rect 564299 312306 564333 312334
rect 564299 312234 564333 312266
rect 564299 312164 564333 312198
rect 564299 312096 564333 312128
rect 564299 312028 564333 312056
rect 564299 311960 564333 311984
rect 564299 311892 564333 311912
rect 564299 311824 564333 311840
rect 564299 311756 564333 311768
rect 564299 311677 564333 311696
rect 564557 312666 564591 312685
rect 564557 312594 564591 312606
rect 564557 312522 564591 312538
rect 564557 312450 564591 312470
rect 564557 312378 564591 312402
rect 564557 312306 564591 312334
rect 564557 312234 564591 312266
rect 564557 312164 564591 312198
rect 564557 312096 564591 312128
rect 564557 312028 564591 312056
rect 564557 311960 564591 311984
rect 564557 311892 564591 311912
rect 564557 311824 564591 311840
rect 564557 311756 564591 311768
rect 564557 311611 564591 311696
rect 564815 312666 564849 312871
rect 564815 312594 564849 312606
rect 564815 312522 564849 312538
rect 564815 312450 564849 312470
rect 564815 312378 564849 312402
rect 564815 312306 564849 312334
rect 564815 312234 564849 312266
rect 564815 312164 564849 312198
rect 564815 312096 564849 312128
rect 564815 312028 564849 312056
rect 564815 311960 564849 311984
rect 564815 311892 564849 311912
rect 564815 311824 564849 311840
rect 564815 311756 564849 311768
rect 564815 311677 564849 311696
rect 565073 312666 565107 312685
rect 565073 312594 565107 312606
rect 565073 312522 565107 312538
rect 565073 312450 565107 312470
rect 565073 312378 565107 312402
rect 565073 312306 565107 312334
rect 565073 312234 565107 312266
rect 565073 312164 565107 312198
rect 565073 312096 565107 312128
rect 565073 312028 565107 312056
rect 565073 311960 565107 311984
rect 565073 311892 565107 311912
rect 565073 311824 565107 311840
rect 565073 311756 565107 311768
rect 565073 311611 565107 311696
rect 565331 312666 565365 312871
rect 565331 312594 565365 312606
rect 565331 312522 565365 312538
rect 565331 312450 565365 312470
rect 565331 312378 565365 312402
rect 565331 312306 565365 312334
rect 565331 312234 565365 312266
rect 565331 312164 565365 312198
rect 565331 312096 565365 312128
rect 565331 312028 565365 312056
rect 565331 311960 565365 311984
rect 565331 311892 565365 311912
rect 565331 311824 565365 311840
rect 565331 311756 565365 311768
rect 565331 311677 565365 311696
rect 565589 312666 565623 312685
rect 565589 312594 565623 312606
rect 565589 312522 565623 312538
rect 565589 312450 565623 312470
rect 565589 312378 565623 312402
rect 565589 312306 565623 312334
rect 565589 312234 565623 312266
rect 565589 312164 565623 312198
rect 565589 312096 565623 312128
rect 565589 312028 565623 312056
rect 565589 311960 565623 311984
rect 565589 311892 565623 311912
rect 565589 311824 565623 311840
rect 565589 311756 565623 311768
rect 565589 311685 565623 311696
rect 565589 311665 565648 311685
rect 565842 311668 566002 311669
rect 565842 311665 565869 311668
rect 565589 311611 565869 311665
rect 560098 311553 560250 311595
rect 560156 311445 560250 311553
rect 560416 311562 565869 311611
rect 565975 311665 566002 311668
rect 565975 311562 566008 311665
rect 574916 311575 574976 312921
rect 575153 312736 575187 312755
rect 575153 312664 575187 312676
rect 575153 312592 575187 312608
rect 575153 312520 575187 312540
rect 575153 312448 575187 312472
rect 575153 312376 575187 312404
rect 575153 312304 575187 312336
rect 575153 312234 575187 312268
rect 575153 312166 575187 312198
rect 575153 312098 575187 312126
rect 575153 312030 575187 312054
rect 575153 311962 575187 311982
rect 575153 311894 575187 311910
rect 575153 311826 575187 311838
rect 575153 311621 575187 311766
rect 575411 312736 575445 312921
rect 575411 312664 575445 312676
rect 575411 312592 575445 312608
rect 575411 312520 575445 312540
rect 575411 312448 575445 312472
rect 575411 312376 575445 312404
rect 575411 312304 575445 312336
rect 575411 312234 575445 312268
rect 575411 312166 575445 312198
rect 575411 312098 575445 312126
rect 575411 312030 575445 312054
rect 575411 311962 575445 311982
rect 575411 311894 575445 311910
rect 575411 311826 575445 311838
rect 575411 311747 575445 311766
rect 575669 312736 575703 312755
rect 575669 312664 575703 312676
rect 575669 312592 575703 312608
rect 575669 312520 575703 312540
rect 575669 312448 575703 312472
rect 575669 312376 575703 312404
rect 575669 312304 575703 312336
rect 575669 312234 575703 312268
rect 575669 312166 575703 312198
rect 575669 312098 575703 312126
rect 575669 312030 575703 312054
rect 575669 311962 575703 311982
rect 575669 311894 575703 311910
rect 575669 311826 575703 311838
rect 575669 311621 575703 311766
rect 575927 312736 575961 312921
rect 575927 312664 575961 312676
rect 575927 312592 575961 312608
rect 575927 312520 575961 312540
rect 575927 312448 575961 312472
rect 575927 312376 575961 312404
rect 575927 312304 575961 312336
rect 575927 312234 575961 312268
rect 575927 312166 575961 312198
rect 575927 312098 575961 312126
rect 575927 312030 575961 312054
rect 575927 311962 575961 311982
rect 575927 311894 575961 311910
rect 575927 311826 575961 311838
rect 575927 311747 575961 311766
rect 576185 312736 576219 312755
rect 576185 312664 576219 312676
rect 576185 312592 576219 312608
rect 576185 312520 576219 312540
rect 576185 312448 576219 312472
rect 576185 312376 576219 312404
rect 576185 312304 576219 312336
rect 576185 312234 576219 312268
rect 576185 312166 576219 312198
rect 576185 312098 576219 312126
rect 576185 312030 576219 312054
rect 576185 311962 576219 311982
rect 576185 311894 576219 311910
rect 576185 311826 576219 311838
rect 576185 311621 576219 311766
rect 576443 312736 576477 312921
rect 576443 312664 576477 312676
rect 576443 312592 576477 312608
rect 576443 312520 576477 312540
rect 576443 312448 576477 312472
rect 576443 312376 576477 312404
rect 576443 312304 576477 312336
rect 576443 312234 576477 312268
rect 576443 312166 576477 312198
rect 576443 312098 576477 312126
rect 576443 312030 576477 312054
rect 576443 311962 576477 311982
rect 576443 311894 576477 311910
rect 576443 311826 576477 311838
rect 576443 311747 576477 311766
rect 576701 312736 576735 312755
rect 576701 312664 576735 312676
rect 576701 312592 576735 312608
rect 576701 312520 576735 312540
rect 576701 312448 576735 312472
rect 576701 312376 576735 312404
rect 576701 312304 576735 312336
rect 576701 312234 576735 312268
rect 576701 312166 576735 312198
rect 576701 312098 576735 312126
rect 576701 312030 576735 312054
rect 576701 311962 576735 311982
rect 576701 311894 576735 311910
rect 576701 311826 576735 311838
rect 576701 311621 576735 311766
rect 576959 312736 576993 312921
rect 576959 312664 576993 312676
rect 576959 312592 576993 312608
rect 576959 312520 576993 312540
rect 576959 312448 576993 312472
rect 576959 312376 576993 312404
rect 576959 312304 576993 312336
rect 576959 312234 576993 312268
rect 576959 312166 576993 312198
rect 576959 312098 576993 312126
rect 576959 312030 576993 312054
rect 576959 311962 576993 311982
rect 576959 311894 576993 311910
rect 576959 311826 576993 311838
rect 576959 311747 576993 311766
rect 577217 312736 577251 312755
rect 577217 312664 577251 312676
rect 577217 312592 577251 312608
rect 577217 312520 577251 312540
rect 577217 312448 577251 312472
rect 577217 312376 577251 312404
rect 577217 312304 577251 312336
rect 577217 312234 577251 312268
rect 577217 312166 577251 312198
rect 577217 312098 577251 312126
rect 577217 312030 577251 312054
rect 577217 311962 577251 311982
rect 577217 311894 577251 311910
rect 577217 311826 577251 311838
rect 577217 311621 577251 311766
rect 577475 312736 577509 312921
rect 577475 312664 577509 312676
rect 577475 312592 577509 312608
rect 577475 312520 577509 312540
rect 577475 312448 577509 312472
rect 577475 312376 577509 312404
rect 577475 312304 577509 312336
rect 577475 312234 577509 312268
rect 577475 312166 577509 312198
rect 577475 312098 577509 312126
rect 577475 312030 577509 312054
rect 577475 311962 577509 311982
rect 577475 311894 577509 311910
rect 577475 311826 577509 311838
rect 577475 311747 577509 311766
rect 577733 312736 577767 312755
rect 577733 312664 577767 312676
rect 577733 312592 577767 312608
rect 577733 312520 577767 312540
rect 577733 312448 577767 312472
rect 577733 312376 577767 312404
rect 577733 312304 577767 312336
rect 577733 312234 577767 312268
rect 577733 312166 577767 312198
rect 577733 312098 577767 312126
rect 577733 312030 577767 312054
rect 577733 311962 577767 311982
rect 577733 311894 577767 311910
rect 577733 311826 577767 311838
rect 577733 311621 577767 311766
rect 577991 312736 578025 312921
rect 577991 312664 578025 312676
rect 577991 312592 578025 312608
rect 577991 312520 578025 312540
rect 577991 312448 578025 312472
rect 577991 312376 578025 312404
rect 577991 312304 578025 312336
rect 577991 312234 578025 312268
rect 577991 312166 578025 312198
rect 577991 312098 578025 312126
rect 577991 312030 578025 312054
rect 577991 311962 578025 311982
rect 577991 311894 578025 311910
rect 577991 311826 578025 311838
rect 577991 311747 578025 311766
rect 578249 312736 578283 312755
rect 578249 312664 578283 312676
rect 578249 312592 578283 312608
rect 578249 312520 578283 312540
rect 578249 312448 578283 312472
rect 578249 312376 578283 312404
rect 578249 312304 578283 312336
rect 578249 312234 578283 312268
rect 578249 312166 578283 312198
rect 578249 312098 578283 312126
rect 578249 312030 578283 312054
rect 578249 311962 578283 311982
rect 578249 311894 578283 311910
rect 578249 311826 578283 311838
rect 578249 311621 578283 311766
rect 578507 312736 578541 312921
rect 578507 312664 578541 312676
rect 578507 312592 578541 312608
rect 578507 312520 578541 312540
rect 578507 312448 578541 312472
rect 578507 312376 578541 312404
rect 578507 312304 578541 312336
rect 578507 312234 578541 312268
rect 578507 312166 578541 312198
rect 578507 312098 578541 312126
rect 578507 312030 578541 312054
rect 578507 311962 578541 311982
rect 578507 311894 578541 311910
rect 578507 311826 578541 311838
rect 578507 311747 578541 311766
rect 578765 312736 578799 312755
rect 578765 312664 578799 312676
rect 578765 312592 578799 312608
rect 578765 312520 578799 312540
rect 578765 312448 578799 312472
rect 578765 312376 578799 312404
rect 578765 312304 578799 312336
rect 578765 312234 578799 312268
rect 578765 312166 578799 312198
rect 578765 312098 578799 312126
rect 578765 312030 578799 312054
rect 578765 311962 578799 311982
rect 578765 311894 578799 311910
rect 578765 311826 578799 311838
rect 578765 311621 578799 311766
rect 579023 312736 579057 312921
rect 579023 312664 579057 312676
rect 579023 312592 579057 312608
rect 579023 312520 579057 312540
rect 579023 312448 579057 312472
rect 579023 312376 579057 312404
rect 579023 312304 579057 312336
rect 579023 312234 579057 312268
rect 579023 312166 579057 312198
rect 579023 312098 579057 312126
rect 579023 312030 579057 312054
rect 579023 311962 579057 311982
rect 579023 311894 579057 311910
rect 579023 311826 579057 311838
rect 579023 311747 579057 311766
rect 579281 312736 579315 312755
rect 579281 312664 579315 312676
rect 579281 312592 579315 312608
rect 579281 312520 579315 312540
rect 579281 312448 579315 312472
rect 579281 312376 579315 312404
rect 579281 312304 579315 312336
rect 579281 312234 579315 312268
rect 579281 312166 579315 312198
rect 579281 312098 579315 312126
rect 579281 312030 579315 312054
rect 579281 311962 579315 311982
rect 579281 311894 579315 311910
rect 579281 311826 579315 311838
rect 579281 311621 579315 311766
rect 579539 312736 579573 312921
rect 579539 312664 579573 312676
rect 579539 312592 579573 312608
rect 579539 312520 579573 312540
rect 579539 312448 579573 312472
rect 579539 312376 579573 312404
rect 579539 312304 579573 312336
rect 579539 312234 579573 312268
rect 579539 312166 579573 312198
rect 579539 312098 579573 312126
rect 579539 312030 579573 312054
rect 579539 311962 579573 311982
rect 579539 311894 579573 311910
rect 579539 311826 579573 311838
rect 579539 311747 579573 311766
rect 579797 312736 579831 312755
rect 579797 312664 579831 312676
rect 579797 312592 579831 312608
rect 579797 312520 579831 312540
rect 579797 312448 579831 312472
rect 579797 312376 579831 312404
rect 579797 312304 579831 312336
rect 579797 312234 579831 312268
rect 579797 312166 579831 312198
rect 579797 312098 579831 312126
rect 579797 312030 579831 312054
rect 579797 311962 579831 311982
rect 579797 311894 579831 311910
rect 579797 311826 579831 311838
rect 579797 311621 579831 311766
rect 580055 312736 580089 312921
rect 580404 312891 580464 312974
rect 580055 312664 580089 312676
rect 580055 312592 580089 312608
rect 580055 312520 580089 312540
rect 580055 312448 580089 312472
rect 580055 312376 580089 312404
rect 580055 312304 580089 312336
rect 580055 312234 580089 312268
rect 580055 312166 580089 312198
rect 580055 312098 580089 312126
rect 580055 312030 580089 312054
rect 580055 311962 580089 311982
rect 580055 311894 580089 311910
rect 580055 311826 580089 311838
rect 580055 311747 580089 311766
rect 580313 312736 580347 312755
rect 580313 312664 580347 312676
rect 580313 312592 580347 312608
rect 580313 312520 580347 312540
rect 580313 312448 580347 312472
rect 580313 312376 580347 312404
rect 580313 312304 580347 312336
rect 580313 312234 580347 312268
rect 580313 312166 580347 312198
rect 580313 312098 580347 312126
rect 580313 312030 580347 312054
rect 580313 311962 580347 311982
rect 580313 311894 580347 311910
rect 580313 311826 580347 311838
rect 580313 311745 580347 311766
rect 580350 311628 580578 311665
rect 580350 311621 580506 311628
rect 560416 311551 566008 311562
rect 574860 311486 574976 311575
rect 575100 311594 580506 311621
rect 580540 311594 580578 311628
rect 575100 311561 580578 311594
rect 574860 311452 574899 311486
rect 574933 311459 574976 311486
rect 574933 311452 580394 311459
rect 574860 311446 580394 311452
rect 560156 311432 565554 311445
rect 560156 311398 560617 311432
rect 560651 311398 560817 311432
rect 560851 311398 561017 311432
rect 561051 311398 561217 311432
rect 561251 311398 561417 311432
rect 561451 311398 561617 311432
rect 561651 311398 561817 311432
rect 561851 311398 562017 311432
rect 562051 311398 562217 311432
rect 562251 311398 562417 311432
rect 562451 311398 562617 311432
rect 562651 311398 562817 311432
rect 562851 311398 563017 311432
rect 563051 311398 563217 311432
rect 563251 311398 563417 311432
rect 563451 311398 563617 311432
rect 563651 311398 563817 311432
rect 563851 311398 564017 311432
rect 564051 311398 564217 311432
rect 564251 311398 564417 311432
rect 564451 311398 564617 311432
rect 564651 311398 564817 311432
rect 564851 311398 565017 311432
rect 565051 311398 565217 311432
rect 565251 311398 565417 311432
rect 565451 311398 565554 311432
rect 560156 311385 565554 311398
rect 565644 311338 565704 311421
rect 574860 311412 575177 311446
rect 575211 311412 575377 311446
rect 575411 311412 575577 311446
rect 575611 311412 575777 311446
rect 575811 311412 575977 311446
rect 576011 311412 576177 311446
rect 576211 311412 576377 311446
rect 576411 311412 576577 311446
rect 576611 311412 576777 311446
rect 576811 311412 576977 311446
rect 577011 311412 577177 311446
rect 577211 311412 577377 311446
rect 577411 311412 577577 311446
rect 577611 311412 577777 311446
rect 577811 311412 577977 311446
rect 578011 311412 578177 311446
rect 578211 311412 578377 311446
rect 578411 311412 578577 311446
rect 578611 311412 578777 311446
rect 578811 311412 578977 311446
rect 579011 311412 579177 311446
rect 579211 311412 579377 311446
rect 579411 311412 579577 311446
rect 579611 311412 579777 311446
rect 579811 311412 579977 311446
rect 580011 311412 580177 311446
rect 580211 311412 580394 311446
rect 574860 311401 580394 311412
rect 574898 311399 580394 311401
rect 561896 311308 562056 311331
rect 561896 311274 561957 311308
rect 561991 311274 562056 311308
rect 561896 311211 562056 311274
rect 563196 311308 563356 311331
rect 563196 311274 563257 311308
rect 563291 311274 563356 311308
rect 563196 311211 563356 311274
rect 564496 311308 564656 311331
rect 564496 311274 564557 311308
rect 564591 311274 564656 311308
rect 564496 311211 564656 311274
rect 565644 311304 565657 311338
rect 565691 311304 565704 311338
rect 565644 311211 565704 311304
rect 575106 311268 580492 311281
rect 575106 311234 575177 311268
rect 575211 311234 575377 311268
rect 575411 311234 575577 311268
rect 575611 311234 575777 311268
rect 575811 311234 575977 311268
rect 576011 311234 576177 311268
rect 576211 311234 576377 311268
rect 576411 311234 576577 311268
rect 576611 311234 576777 311268
rect 576811 311234 576977 311268
rect 577011 311234 577177 311268
rect 577211 311234 577377 311268
rect 577411 311234 577577 311268
rect 577611 311234 577777 311268
rect 577811 311234 577977 311268
rect 578011 311234 578177 311268
rect 578211 311234 578377 311268
rect 578411 311234 578577 311268
rect 578611 311234 578777 311268
rect 578811 311234 578977 311268
rect 579011 311234 579177 311268
rect 579211 311234 579377 311268
rect 579411 311234 579577 311268
rect 579611 311234 579777 311268
rect 579811 311234 579977 311268
rect 580011 311234 580177 311268
rect 580211 311234 580492 311268
rect 575106 311221 580492 311234
rect 560418 311198 565732 311211
rect 560418 311164 560617 311198
rect 560651 311164 560817 311198
rect 560851 311164 561017 311198
rect 561051 311164 561217 311198
rect 561251 311164 561417 311198
rect 561451 311164 561617 311198
rect 561651 311164 561817 311198
rect 561851 311164 562017 311198
rect 562051 311164 562217 311198
rect 562251 311164 562417 311198
rect 562451 311164 562617 311198
rect 562651 311164 562817 311198
rect 562851 311164 563017 311198
rect 563051 311164 563217 311198
rect 563251 311164 563417 311198
rect 563451 311164 563617 311198
rect 563651 311164 563817 311198
rect 563851 311164 564017 311198
rect 564051 311164 564217 311198
rect 564251 311164 564417 311198
rect 564451 311164 564617 311198
rect 564651 311164 564817 311198
rect 564851 311164 565017 311198
rect 565051 311164 565217 311198
rect 565251 311164 565417 311198
rect 565451 311164 565732 311198
rect 560418 311151 565732 311164
<< viali >>
rect 560863 493812 560897 493846
rect 561063 493812 561097 493846
rect 561263 493812 561297 493846
rect 561463 493812 561497 493846
rect 561663 493812 561697 493846
rect 561863 493812 561897 493846
rect 562063 493812 562097 493846
rect 562263 493812 562297 493846
rect 562463 493812 562497 493846
rect 562663 493812 562697 493846
rect 562863 493812 562897 493846
rect 563063 493812 563097 493846
rect 563263 493812 563297 493846
rect 563463 493812 563497 493846
rect 563663 493812 563697 493846
rect 563863 493812 563897 493846
rect 564063 493812 564097 493846
rect 564263 493812 564297 493846
rect 564463 493812 564497 493846
rect 564663 493812 564697 493846
rect 564863 493812 564897 493846
rect 565063 493812 565097 493846
rect 565263 493812 565297 493846
rect 565463 493812 565497 493846
rect 565663 493812 565697 493846
rect 560367 492363 560473 492469
rect 560675 493408 560709 493434
rect 560675 493400 560709 493408
rect 560675 493340 560709 493362
rect 560675 493328 560709 493340
rect 560675 493272 560709 493290
rect 560675 493256 560709 493272
rect 560675 493204 560709 493218
rect 560675 493184 560709 493204
rect 560675 493136 560709 493146
rect 560675 493112 560709 493136
rect 560675 493068 560709 493074
rect 560675 493040 560709 493068
rect 560675 493000 560709 493002
rect 560675 492968 560709 493000
rect 560675 492898 560709 492930
rect 560675 492896 560709 492898
rect 560675 492830 560709 492858
rect 560675 492824 560709 492830
rect 560675 492762 560709 492786
rect 560675 492752 560709 492762
rect 560675 492694 560709 492714
rect 560675 492680 560709 492694
rect 560675 492626 560709 492642
rect 560675 492608 560709 492626
rect 560675 492558 560709 492570
rect 560675 492536 560709 492558
rect 560675 492490 560709 492498
rect 560675 492464 560709 492490
rect 560933 493408 560967 493434
rect 560933 493400 560967 493408
rect 560933 493340 560967 493362
rect 560933 493328 560967 493340
rect 560933 493272 560967 493290
rect 560933 493256 560967 493272
rect 560933 493204 560967 493218
rect 560933 493184 560967 493204
rect 560933 493136 560967 493146
rect 560933 493112 560967 493136
rect 560933 493068 560967 493074
rect 560933 493040 560967 493068
rect 560933 493000 560967 493002
rect 560933 492968 560967 493000
rect 560933 492898 560967 492930
rect 560933 492896 560967 492898
rect 560933 492830 560967 492858
rect 560933 492824 560967 492830
rect 560933 492762 560967 492786
rect 560933 492752 560967 492762
rect 560933 492694 560967 492714
rect 560933 492680 560967 492694
rect 560933 492626 560967 492642
rect 560933 492608 560967 492626
rect 560933 492558 560967 492570
rect 560933 492536 560967 492558
rect 560933 492490 560967 492498
rect 560933 492464 560967 492490
rect 561191 493408 561225 493434
rect 561191 493400 561225 493408
rect 561191 493340 561225 493362
rect 561191 493328 561225 493340
rect 561191 493272 561225 493290
rect 561191 493256 561225 493272
rect 561191 493204 561225 493218
rect 561191 493184 561225 493204
rect 561191 493136 561225 493146
rect 561191 493112 561225 493136
rect 561191 493068 561225 493074
rect 561191 493040 561225 493068
rect 561191 493000 561225 493002
rect 561191 492968 561225 493000
rect 561191 492898 561225 492930
rect 561191 492896 561225 492898
rect 561191 492830 561225 492858
rect 561191 492824 561225 492830
rect 561191 492762 561225 492786
rect 561191 492752 561225 492762
rect 561191 492694 561225 492714
rect 561191 492680 561225 492694
rect 561191 492626 561225 492642
rect 561191 492608 561225 492626
rect 561191 492558 561225 492570
rect 561191 492536 561225 492558
rect 561191 492490 561225 492498
rect 561191 492464 561225 492490
rect 561449 493408 561483 493434
rect 561449 493400 561483 493408
rect 561449 493340 561483 493362
rect 561449 493328 561483 493340
rect 561449 493272 561483 493290
rect 561449 493256 561483 493272
rect 561449 493204 561483 493218
rect 561449 493184 561483 493204
rect 561449 493136 561483 493146
rect 561449 493112 561483 493136
rect 561449 493068 561483 493074
rect 561449 493040 561483 493068
rect 561449 493000 561483 493002
rect 561449 492968 561483 493000
rect 561449 492898 561483 492930
rect 561449 492896 561483 492898
rect 561449 492830 561483 492858
rect 561449 492824 561483 492830
rect 561449 492762 561483 492786
rect 561449 492752 561483 492762
rect 561449 492694 561483 492714
rect 561449 492680 561483 492694
rect 561449 492626 561483 492642
rect 561449 492608 561483 492626
rect 561449 492558 561483 492570
rect 561449 492536 561483 492558
rect 561449 492490 561483 492498
rect 561449 492464 561483 492490
rect 561707 493408 561741 493434
rect 561707 493400 561741 493408
rect 561707 493340 561741 493362
rect 561707 493328 561741 493340
rect 561707 493272 561741 493290
rect 561707 493256 561741 493272
rect 561707 493204 561741 493218
rect 561707 493184 561741 493204
rect 561707 493136 561741 493146
rect 561707 493112 561741 493136
rect 561707 493068 561741 493074
rect 561707 493040 561741 493068
rect 561707 493000 561741 493002
rect 561707 492968 561741 493000
rect 561707 492898 561741 492930
rect 561707 492896 561741 492898
rect 561707 492830 561741 492858
rect 561707 492824 561741 492830
rect 561707 492762 561741 492786
rect 561707 492752 561741 492762
rect 561707 492694 561741 492714
rect 561707 492680 561741 492694
rect 561707 492626 561741 492642
rect 561707 492608 561741 492626
rect 561707 492558 561741 492570
rect 561707 492536 561741 492558
rect 561707 492490 561741 492498
rect 561707 492464 561741 492490
rect 561965 493408 561999 493434
rect 561965 493400 561999 493408
rect 561965 493340 561999 493362
rect 561965 493328 561999 493340
rect 561965 493272 561999 493290
rect 561965 493256 561999 493272
rect 561965 493204 561999 493218
rect 561965 493184 561999 493204
rect 561965 493136 561999 493146
rect 561965 493112 561999 493136
rect 561965 493068 561999 493074
rect 561965 493040 561999 493068
rect 561965 493000 561999 493002
rect 561965 492968 561999 493000
rect 561965 492898 561999 492930
rect 561965 492896 561999 492898
rect 561965 492830 561999 492858
rect 561965 492824 561999 492830
rect 561965 492762 561999 492786
rect 561965 492752 561999 492762
rect 561965 492694 561999 492714
rect 561965 492680 561999 492694
rect 561965 492626 561999 492642
rect 561965 492608 561999 492626
rect 561965 492558 561999 492570
rect 561965 492536 561999 492558
rect 561965 492490 561999 492498
rect 561965 492464 561999 492490
rect 562223 493408 562257 493434
rect 562223 493400 562257 493408
rect 562223 493340 562257 493362
rect 562223 493328 562257 493340
rect 562223 493272 562257 493290
rect 562223 493256 562257 493272
rect 562223 493204 562257 493218
rect 562223 493184 562257 493204
rect 562223 493136 562257 493146
rect 562223 493112 562257 493136
rect 562223 493068 562257 493074
rect 562223 493040 562257 493068
rect 562223 493000 562257 493002
rect 562223 492968 562257 493000
rect 562223 492898 562257 492930
rect 562223 492896 562257 492898
rect 562223 492830 562257 492858
rect 562223 492824 562257 492830
rect 562223 492762 562257 492786
rect 562223 492752 562257 492762
rect 562223 492694 562257 492714
rect 562223 492680 562257 492694
rect 562223 492626 562257 492642
rect 562223 492608 562257 492626
rect 562223 492558 562257 492570
rect 562223 492536 562257 492558
rect 562223 492490 562257 492498
rect 562223 492464 562257 492490
rect 562481 493408 562515 493434
rect 562481 493400 562515 493408
rect 562481 493340 562515 493362
rect 562481 493328 562515 493340
rect 562481 493272 562515 493290
rect 562481 493256 562515 493272
rect 562481 493204 562515 493218
rect 562481 493184 562515 493204
rect 562481 493136 562515 493146
rect 562481 493112 562515 493136
rect 562481 493068 562515 493074
rect 562481 493040 562515 493068
rect 562481 493000 562515 493002
rect 562481 492968 562515 493000
rect 562481 492898 562515 492930
rect 562481 492896 562515 492898
rect 562481 492830 562515 492858
rect 562481 492824 562515 492830
rect 562481 492762 562515 492786
rect 562481 492752 562515 492762
rect 562481 492694 562515 492714
rect 562481 492680 562515 492694
rect 562481 492626 562515 492642
rect 562481 492608 562515 492626
rect 562481 492558 562515 492570
rect 562481 492536 562515 492558
rect 562481 492490 562515 492498
rect 562481 492464 562515 492490
rect 562739 493408 562773 493434
rect 562739 493400 562773 493408
rect 562739 493340 562773 493362
rect 562739 493328 562773 493340
rect 562739 493272 562773 493290
rect 562739 493256 562773 493272
rect 562739 493204 562773 493218
rect 562739 493184 562773 493204
rect 562739 493136 562773 493146
rect 562739 493112 562773 493136
rect 562739 493068 562773 493074
rect 562739 493040 562773 493068
rect 562739 493000 562773 493002
rect 562739 492968 562773 493000
rect 562739 492898 562773 492930
rect 562739 492896 562773 492898
rect 562739 492830 562773 492858
rect 562739 492824 562773 492830
rect 562739 492762 562773 492786
rect 562739 492752 562773 492762
rect 562739 492694 562773 492714
rect 562739 492680 562773 492694
rect 562739 492626 562773 492642
rect 562739 492608 562773 492626
rect 562739 492558 562773 492570
rect 562739 492536 562773 492558
rect 562739 492490 562773 492498
rect 562739 492464 562773 492490
rect 562997 493408 563031 493434
rect 562997 493400 563031 493408
rect 562997 493340 563031 493362
rect 562997 493328 563031 493340
rect 562997 493272 563031 493290
rect 562997 493256 563031 493272
rect 562997 493204 563031 493218
rect 562997 493184 563031 493204
rect 562997 493136 563031 493146
rect 562997 493112 563031 493136
rect 562997 493068 563031 493074
rect 562997 493040 563031 493068
rect 562997 493000 563031 493002
rect 562997 492968 563031 493000
rect 562997 492898 563031 492930
rect 562997 492896 563031 492898
rect 562997 492830 563031 492858
rect 562997 492824 563031 492830
rect 562997 492762 563031 492786
rect 562997 492752 563031 492762
rect 562997 492694 563031 492714
rect 562997 492680 563031 492694
rect 562997 492626 563031 492642
rect 562997 492608 563031 492626
rect 562997 492558 563031 492570
rect 562997 492536 563031 492558
rect 562997 492490 563031 492498
rect 562997 492464 563031 492490
rect 563255 493408 563289 493434
rect 563255 493400 563289 493408
rect 563255 493340 563289 493362
rect 563255 493328 563289 493340
rect 563255 493272 563289 493290
rect 563255 493256 563289 493272
rect 563255 493204 563289 493218
rect 563255 493184 563289 493204
rect 563255 493136 563289 493146
rect 563255 493112 563289 493136
rect 563255 493068 563289 493074
rect 563255 493040 563289 493068
rect 563255 493000 563289 493002
rect 563255 492968 563289 493000
rect 563255 492898 563289 492930
rect 563255 492896 563289 492898
rect 563255 492830 563289 492858
rect 563255 492824 563289 492830
rect 563255 492762 563289 492786
rect 563255 492752 563289 492762
rect 563255 492694 563289 492714
rect 563255 492680 563289 492694
rect 563255 492626 563289 492642
rect 563255 492608 563289 492626
rect 563255 492558 563289 492570
rect 563255 492536 563289 492558
rect 563255 492490 563289 492498
rect 563255 492464 563289 492490
rect 563513 493408 563547 493434
rect 563513 493400 563547 493408
rect 563513 493340 563547 493362
rect 563513 493328 563547 493340
rect 563513 493272 563547 493290
rect 563513 493256 563547 493272
rect 563513 493204 563547 493218
rect 563513 493184 563547 493204
rect 563513 493136 563547 493146
rect 563513 493112 563547 493136
rect 563513 493068 563547 493074
rect 563513 493040 563547 493068
rect 563513 493000 563547 493002
rect 563513 492968 563547 493000
rect 563513 492898 563547 492930
rect 563513 492896 563547 492898
rect 563513 492830 563547 492858
rect 563513 492824 563547 492830
rect 563513 492762 563547 492786
rect 563513 492752 563547 492762
rect 563513 492694 563547 492714
rect 563513 492680 563547 492694
rect 563513 492626 563547 492642
rect 563513 492608 563547 492626
rect 563513 492558 563547 492570
rect 563513 492536 563547 492558
rect 563513 492490 563547 492498
rect 563513 492464 563547 492490
rect 563771 493408 563805 493434
rect 563771 493400 563805 493408
rect 563771 493340 563805 493362
rect 563771 493328 563805 493340
rect 563771 493272 563805 493290
rect 563771 493256 563805 493272
rect 563771 493204 563805 493218
rect 563771 493184 563805 493204
rect 563771 493136 563805 493146
rect 563771 493112 563805 493136
rect 563771 493068 563805 493074
rect 563771 493040 563805 493068
rect 563771 493000 563805 493002
rect 563771 492968 563805 493000
rect 563771 492898 563805 492930
rect 563771 492896 563805 492898
rect 563771 492830 563805 492858
rect 563771 492824 563805 492830
rect 563771 492762 563805 492786
rect 563771 492752 563805 492762
rect 563771 492694 563805 492714
rect 563771 492680 563805 492694
rect 563771 492626 563805 492642
rect 563771 492608 563805 492626
rect 563771 492558 563805 492570
rect 563771 492536 563805 492558
rect 563771 492490 563805 492498
rect 563771 492464 563805 492490
rect 564029 493408 564063 493434
rect 564029 493400 564063 493408
rect 564029 493340 564063 493362
rect 564029 493328 564063 493340
rect 564029 493272 564063 493290
rect 564029 493256 564063 493272
rect 564029 493204 564063 493218
rect 564029 493184 564063 493204
rect 564029 493136 564063 493146
rect 564029 493112 564063 493136
rect 564029 493068 564063 493074
rect 564029 493040 564063 493068
rect 564029 493000 564063 493002
rect 564029 492968 564063 493000
rect 564029 492898 564063 492930
rect 564029 492896 564063 492898
rect 564029 492830 564063 492858
rect 564029 492824 564063 492830
rect 564029 492762 564063 492786
rect 564029 492752 564063 492762
rect 564029 492694 564063 492714
rect 564029 492680 564063 492694
rect 564029 492626 564063 492642
rect 564029 492608 564063 492626
rect 564029 492558 564063 492570
rect 564029 492536 564063 492558
rect 564029 492490 564063 492498
rect 564029 492464 564063 492490
rect 564287 493408 564321 493434
rect 564287 493400 564321 493408
rect 564287 493340 564321 493362
rect 564287 493328 564321 493340
rect 564287 493272 564321 493290
rect 564287 493256 564321 493272
rect 564287 493204 564321 493218
rect 564287 493184 564321 493204
rect 564287 493136 564321 493146
rect 564287 493112 564321 493136
rect 564287 493068 564321 493074
rect 564287 493040 564321 493068
rect 564287 493000 564321 493002
rect 564287 492968 564321 493000
rect 564287 492898 564321 492930
rect 564287 492896 564321 492898
rect 564287 492830 564321 492858
rect 564287 492824 564321 492830
rect 564287 492762 564321 492786
rect 564287 492752 564321 492762
rect 564287 492694 564321 492714
rect 564287 492680 564321 492694
rect 564287 492626 564321 492642
rect 564287 492608 564321 492626
rect 564287 492558 564321 492570
rect 564287 492536 564321 492558
rect 564287 492490 564321 492498
rect 564287 492464 564321 492490
rect 564545 493408 564579 493434
rect 564545 493400 564579 493408
rect 564545 493340 564579 493362
rect 564545 493328 564579 493340
rect 564545 493272 564579 493290
rect 564545 493256 564579 493272
rect 564545 493204 564579 493218
rect 564545 493184 564579 493204
rect 564545 493136 564579 493146
rect 564545 493112 564579 493136
rect 564545 493068 564579 493074
rect 564545 493040 564579 493068
rect 564545 493000 564579 493002
rect 564545 492968 564579 493000
rect 564545 492898 564579 492930
rect 564545 492896 564579 492898
rect 564545 492830 564579 492858
rect 564545 492824 564579 492830
rect 564545 492762 564579 492786
rect 564545 492752 564579 492762
rect 564545 492694 564579 492714
rect 564545 492680 564579 492694
rect 564545 492626 564579 492642
rect 564545 492608 564579 492626
rect 564545 492558 564579 492570
rect 564545 492536 564579 492558
rect 564545 492490 564579 492498
rect 564545 492464 564579 492490
rect 564803 493408 564837 493434
rect 564803 493400 564837 493408
rect 564803 493340 564837 493362
rect 564803 493328 564837 493340
rect 564803 493272 564837 493290
rect 564803 493256 564837 493272
rect 564803 493204 564837 493218
rect 564803 493184 564837 493204
rect 564803 493136 564837 493146
rect 564803 493112 564837 493136
rect 564803 493068 564837 493074
rect 564803 493040 564837 493068
rect 564803 493000 564837 493002
rect 564803 492968 564837 493000
rect 564803 492898 564837 492930
rect 564803 492896 564837 492898
rect 564803 492830 564837 492858
rect 564803 492824 564837 492830
rect 564803 492762 564837 492786
rect 564803 492752 564837 492762
rect 564803 492694 564837 492714
rect 564803 492680 564837 492694
rect 564803 492626 564837 492642
rect 564803 492608 564837 492626
rect 564803 492558 564837 492570
rect 564803 492536 564837 492558
rect 564803 492490 564837 492498
rect 564803 492464 564837 492490
rect 565061 493408 565095 493434
rect 565061 493400 565095 493408
rect 565061 493340 565095 493362
rect 565061 493328 565095 493340
rect 565061 493272 565095 493290
rect 565061 493256 565095 493272
rect 565061 493204 565095 493218
rect 565061 493184 565095 493204
rect 565061 493136 565095 493146
rect 565061 493112 565095 493136
rect 565061 493068 565095 493074
rect 565061 493040 565095 493068
rect 565061 493000 565095 493002
rect 565061 492968 565095 493000
rect 565061 492898 565095 492930
rect 565061 492896 565095 492898
rect 565061 492830 565095 492858
rect 565061 492824 565095 492830
rect 565061 492762 565095 492786
rect 565061 492752 565095 492762
rect 565061 492694 565095 492714
rect 565061 492680 565095 492694
rect 565061 492626 565095 492642
rect 565061 492608 565095 492626
rect 565061 492558 565095 492570
rect 565061 492536 565095 492558
rect 565061 492490 565095 492498
rect 565061 492464 565095 492490
rect 565319 493408 565353 493434
rect 565319 493400 565353 493408
rect 565319 493340 565353 493362
rect 565319 493328 565353 493340
rect 565319 493272 565353 493290
rect 565319 493256 565353 493272
rect 565319 493204 565353 493218
rect 565319 493184 565353 493204
rect 565319 493136 565353 493146
rect 565319 493112 565353 493136
rect 565319 493068 565353 493074
rect 565319 493040 565353 493068
rect 565319 493000 565353 493002
rect 565319 492968 565353 493000
rect 565319 492898 565353 492930
rect 565319 492896 565353 492898
rect 565319 492830 565353 492858
rect 565319 492824 565353 492830
rect 565319 492762 565353 492786
rect 565319 492752 565353 492762
rect 565319 492694 565353 492714
rect 565319 492680 565353 492694
rect 565319 492626 565353 492642
rect 565319 492608 565353 492626
rect 565319 492558 565353 492570
rect 565319 492536 565353 492558
rect 565319 492490 565353 492498
rect 565319 492464 565353 492490
rect 575255 493586 575289 493620
rect 575455 493586 575489 493620
rect 575655 493586 575689 493620
rect 575855 493586 575889 493620
rect 576055 493586 576089 493620
rect 576255 493586 576289 493620
rect 576455 493586 576489 493620
rect 576655 493586 576689 493620
rect 576855 493586 576889 493620
rect 577055 493586 577089 493620
rect 577255 493586 577289 493620
rect 577455 493586 577489 493620
rect 577655 493586 577689 493620
rect 577855 493586 577889 493620
rect 578055 493586 578089 493620
rect 578255 493586 578289 493620
rect 578455 493586 578489 493620
rect 578655 493586 578689 493620
rect 578855 493586 578889 493620
rect 579055 493586 579089 493620
rect 579255 493586 579289 493620
rect 579455 493586 579489 493620
rect 579655 493586 579689 493620
rect 579855 493586 579889 493620
rect 580055 493586 580089 493620
rect 580255 493586 580289 493620
rect 565577 493408 565611 493434
rect 565577 493400 565611 493408
rect 565577 493340 565611 493362
rect 565577 493328 565611 493340
rect 565577 493272 565611 493290
rect 565577 493256 565611 493272
rect 565577 493204 565611 493218
rect 565577 493184 565611 493204
rect 565577 493136 565611 493146
rect 565577 493112 565611 493136
rect 565577 493068 565611 493074
rect 565577 493040 565611 493068
rect 565577 493000 565611 493002
rect 565577 492968 565611 493000
rect 565577 492898 565611 492930
rect 565577 492896 565611 492898
rect 565577 492830 565611 492858
rect 565577 492824 565611 492830
rect 565577 492762 565611 492786
rect 565577 492752 565611 492762
rect 565577 492694 565611 492714
rect 565577 492680 565611 492694
rect 565577 492626 565611 492642
rect 565577 492608 565611 492626
rect 565577 492558 565611 492570
rect 565577 492536 565611 492558
rect 565577 492490 565611 492498
rect 565577 492464 565611 492490
rect 565835 493408 565869 493434
rect 565835 493400 565869 493408
rect 565835 493340 565869 493362
rect 565835 493328 565869 493340
rect 565835 493272 565869 493290
rect 565835 493256 565869 493272
rect 565835 493204 565869 493218
rect 565835 493184 565869 493204
rect 565835 493136 565869 493146
rect 565835 493112 565869 493136
rect 565835 493068 565869 493074
rect 565835 493040 565869 493068
rect 565835 493000 565869 493002
rect 565835 492968 565869 493000
rect 565835 492898 565869 492930
rect 565835 492896 565869 492898
rect 565835 492830 565869 492858
rect 565835 492824 565869 492830
rect 565835 492762 565869 492786
rect 565835 492752 565869 492762
rect 565835 492694 565869 492714
rect 565835 492680 565869 492694
rect 565835 492626 565869 492642
rect 565835 492608 565869 492626
rect 565835 492558 565869 492570
rect 565835 492536 565869 492558
rect 565835 492490 565869 492498
rect 565835 492464 565869 492490
rect 566115 492330 566221 492436
rect 575231 493182 575265 493208
rect 575231 493174 575265 493182
rect 575231 493114 575265 493136
rect 575231 493102 575265 493114
rect 575231 493046 575265 493064
rect 575231 493030 575265 493046
rect 575231 492978 575265 492992
rect 575231 492958 575265 492978
rect 575231 492910 575265 492920
rect 575231 492886 575265 492910
rect 575231 492842 575265 492848
rect 575231 492814 575265 492842
rect 575231 492774 575265 492776
rect 575231 492742 575265 492774
rect 575231 492672 575265 492704
rect 575231 492670 575265 492672
rect 575231 492604 575265 492632
rect 575231 492598 575265 492604
rect 575231 492536 575265 492560
rect 575231 492526 575265 492536
rect 575231 492468 575265 492488
rect 575231 492454 575265 492468
rect 575231 492400 575265 492416
rect 575231 492382 575265 492400
rect 575231 492332 575265 492344
rect 575231 492310 575265 492332
rect 575231 492264 575265 492272
rect 575231 492238 575265 492264
rect 575489 493182 575523 493208
rect 575489 493174 575523 493182
rect 575489 493114 575523 493136
rect 575489 493102 575523 493114
rect 575489 493046 575523 493064
rect 575489 493030 575523 493046
rect 575489 492978 575523 492992
rect 575489 492958 575523 492978
rect 575489 492910 575523 492920
rect 575489 492886 575523 492910
rect 575489 492842 575523 492848
rect 575489 492814 575523 492842
rect 575489 492774 575523 492776
rect 575489 492742 575523 492774
rect 575489 492672 575523 492704
rect 575489 492670 575523 492672
rect 575489 492604 575523 492632
rect 575489 492598 575523 492604
rect 575489 492536 575523 492560
rect 575489 492526 575523 492536
rect 575489 492468 575523 492488
rect 575489 492454 575523 492468
rect 575489 492400 575523 492416
rect 575489 492382 575523 492400
rect 575489 492332 575523 492344
rect 575489 492310 575523 492332
rect 575489 492264 575523 492272
rect 575489 492238 575523 492264
rect 575747 493182 575781 493208
rect 575747 493174 575781 493182
rect 575747 493114 575781 493136
rect 575747 493102 575781 493114
rect 575747 493046 575781 493064
rect 575747 493030 575781 493046
rect 575747 492978 575781 492992
rect 575747 492958 575781 492978
rect 575747 492910 575781 492920
rect 575747 492886 575781 492910
rect 575747 492842 575781 492848
rect 575747 492814 575781 492842
rect 575747 492774 575781 492776
rect 575747 492742 575781 492774
rect 575747 492672 575781 492704
rect 575747 492670 575781 492672
rect 575747 492604 575781 492632
rect 575747 492598 575781 492604
rect 575747 492536 575781 492560
rect 575747 492526 575781 492536
rect 575747 492468 575781 492488
rect 575747 492454 575781 492468
rect 575747 492400 575781 492416
rect 575747 492382 575781 492400
rect 575747 492332 575781 492344
rect 575747 492310 575781 492332
rect 575747 492264 575781 492272
rect 575747 492238 575781 492264
rect 576005 493182 576039 493208
rect 576005 493174 576039 493182
rect 576005 493114 576039 493136
rect 576005 493102 576039 493114
rect 576005 493046 576039 493064
rect 576005 493030 576039 493046
rect 576005 492978 576039 492992
rect 576005 492958 576039 492978
rect 576005 492910 576039 492920
rect 576005 492886 576039 492910
rect 576005 492842 576039 492848
rect 576005 492814 576039 492842
rect 576005 492774 576039 492776
rect 576005 492742 576039 492774
rect 576005 492672 576039 492704
rect 576005 492670 576039 492672
rect 576005 492604 576039 492632
rect 576005 492598 576039 492604
rect 576005 492536 576039 492560
rect 576005 492526 576039 492536
rect 576005 492468 576039 492488
rect 576005 492454 576039 492468
rect 576005 492400 576039 492416
rect 576005 492382 576039 492400
rect 576005 492332 576039 492344
rect 576005 492310 576039 492332
rect 576005 492264 576039 492272
rect 576005 492238 576039 492264
rect 576263 493182 576297 493208
rect 576263 493174 576297 493182
rect 576263 493114 576297 493136
rect 576263 493102 576297 493114
rect 576263 493046 576297 493064
rect 576263 493030 576297 493046
rect 576263 492978 576297 492992
rect 576263 492958 576297 492978
rect 576263 492910 576297 492920
rect 576263 492886 576297 492910
rect 576263 492842 576297 492848
rect 576263 492814 576297 492842
rect 576263 492774 576297 492776
rect 576263 492742 576297 492774
rect 576263 492672 576297 492704
rect 576263 492670 576297 492672
rect 576263 492604 576297 492632
rect 576263 492598 576297 492604
rect 576263 492536 576297 492560
rect 576263 492526 576297 492536
rect 576263 492468 576297 492488
rect 576263 492454 576297 492468
rect 576263 492400 576297 492416
rect 576263 492382 576297 492400
rect 576263 492332 576297 492344
rect 576263 492310 576297 492332
rect 576263 492264 576297 492272
rect 576263 492238 576297 492264
rect 576521 493182 576555 493208
rect 576521 493174 576555 493182
rect 576521 493114 576555 493136
rect 576521 493102 576555 493114
rect 576521 493046 576555 493064
rect 576521 493030 576555 493046
rect 576521 492978 576555 492992
rect 576521 492958 576555 492978
rect 576521 492910 576555 492920
rect 576521 492886 576555 492910
rect 576521 492842 576555 492848
rect 576521 492814 576555 492842
rect 576521 492774 576555 492776
rect 576521 492742 576555 492774
rect 576521 492672 576555 492704
rect 576521 492670 576555 492672
rect 576521 492604 576555 492632
rect 576521 492598 576555 492604
rect 576521 492536 576555 492560
rect 576521 492526 576555 492536
rect 576521 492468 576555 492488
rect 576521 492454 576555 492468
rect 576521 492400 576555 492416
rect 576521 492382 576555 492400
rect 576521 492332 576555 492344
rect 576521 492310 576555 492332
rect 576521 492264 576555 492272
rect 576521 492238 576555 492264
rect 576779 493182 576813 493208
rect 576779 493174 576813 493182
rect 576779 493114 576813 493136
rect 576779 493102 576813 493114
rect 576779 493046 576813 493064
rect 576779 493030 576813 493046
rect 576779 492978 576813 492992
rect 576779 492958 576813 492978
rect 576779 492910 576813 492920
rect 576779 492886 576813 492910
rect 576779 492842 576813 492848
rect 576779 492814 576813 492842
rect 576779 492774 576813 492776
rect 576779 492742 576813 492774
rect 576779 492672 576813 492704
rect 576779 492670 576813 492672
rect 576779 492604 576813 492632
rect 576779 492598 576813 492604
rect 576779 492536 576813 492560
rect 576779 492526 576813 492536
rect 576779 492468 576813 492488
rect 576779 492454 576813 492468
rect 576779 492400 576813 492416
rect 576779 492382 576813 492400
rect 576779 492332 576813 492344
rect 576779 492310 576813 492332
rect 576779 492264 576813 492272
rect 576779 492238 576813 492264
rect 577037 493182 577071 493208
rect 577037 493174 577071 493182
rect 577037 493114 577071 493136
rect 577037 493102 577071 493114
rect 577037 493046 577071 493064
rect 577037 493030 577071 493046
rect 577037 492978 577071 492992
rect 577037 492958 577071 492978
rect 577037 492910 577071 492920
rect 577037 492886 577071 492910
rect 577037 492842 577071 492848
rect 577037 492814 577071 492842
rect 577037 492774 577071 492776
rect 577037 492742 577071 492774
rect 577037 492672 577071 492704
rect 577037 492670 577071 492672
rect 577037 492604 577071 492632
rect 577037 492598 577071 492604
rect 577037 492536 577071 492560
rect 577037 492526 577071 492536
rect 577037 492468 577071 492488
rect 577037 492454 577071 492468
rect 577037 492400 577071 492416
rect 577037 492382 577071 492400
rect 577037 492332 577071 492344
rect 577037 492310 577071 492332
rect 577037 492264 577071 492272
rect 577037 492238 577071 492264
rect 577295 493182 577329 493208
rect 577295 493174 577329 493182
rect 577295 493114 577329 493136
rect 577295 493102 577329 493114
rect 577295 493046 577329 493064
rect 577295 493030 577329 493046
rect 577295 492978 577329 492992
rect 577295 492958 577329 492978
rect 577295 492910 577329 492920
rect 577295 492886 577329 492910
rect 577295 492842 577329 492848
rect 577295 492814 577329 492842
rect 577295 492774 577329 492776
rect 577295 492742 577329 492774
rect 577295 492672 577329 492704
rect 577295 492670 577329 492672
rect 577295 492604 577329 492632
rect 577295 492598 577329 492604
rect 577295 492536 577329 492560
rect 577295 492526 577329 492536
rect 577295 492468 577329 492488
rect 577295 492454 577329 492468
rect 577295 492400 577329 492416
rect 577295 492382 577329 492400
rect 577295 492332 577329 492344
rect 577295 492310 577329 492332
rect 577295 492264 577329 492272
rect 577295 492238 577329 492264
rect 577553 493182 577587 493208
rect 577553 493174 577587 493182
rect 577553 493114 577587 493136
rect 577553 493102 577587 493114
rect 577553 493046 577587 493064
rect 577553 493030 577587 493046
rect 577553 492978 577587 492992
rect 577553 492958 577587 492978
rect 577553 492910 577587 492920
rect 577553 492886 577587 492910
rect 577553 492842 577587 492848
rect 577553 492814 577587 492842
rect 577553 492774 577587 492776
rect 577553 492742 577587 492774
rect 577553 492672 577587 492704
rect 577553 492670 577587 492672
rect 577553 492604 577587 492632
rect 577553 492598 577587 492604
rect 577553 492536 577587 492560
rect 577553 492526 577587 492536
rect 577553 492468 577587 492488
rect 577553 492454 577587 492468
rect 577553 492400 577587 492416
rect 577553 492382 577587 492400
rect 577553 492332 577587 492344
rect 577553 492310 577587 492332
rect 577553 492264 577587 492272
rect 577553 492238 577587 492264
rect 577811 493182 577845 493208
rect 577811 493174 577845 493182
rect 577811 493114 577845 493136
rect 577811 493102 577845 493114
rect 577811 493046 577845 493064
rect 577811 493030 577845 493046
rect 577811 492978 577845 492992
rect 577811 492958 577845 492978
rect 577811 492910 577845 492920
rect 577811 492886 577845 492910
rect 577811 492842 577845 492848
rect 577811 492814 577845 492842
rect 577811 492774 577845 492776
rect 577811 492742 577845 492774
rect 577811 492672 577845 492704
rect 577811 492670 577845 492672
rect 577811 492604 577845 492632
rect 577811 492598 577845 492604
rect 577811 492536 577845 492560
rect 577811 492526 577845 492536
rect 577811 492468 577845 492488
rect 577811 492454 577845 492468
rect 577811 492400 577845 492416
rect 577811 492382 577845 492400
rect 577811 492332 577845 492344
rect 577811 492310 577845 492332
rect 577811 492264 577845 492272
rect 577811 492238 577845 492264
rect 578069 493182 578103 493208
rect 578069 493174 578103 493182
rect 578069 493114 578103 493136
rect 578069 493102 578103 493114
rect 578069 493046 578103 493064
rect 578069 493030 578103 493046
rect 578069 492978 578103 492992
rect 578069 492958 578103 492978
rect 578069 492910 578103 492920
rect 578069 492886 578103 492910
rect 578069 492842 578103 492848
rect 578069 492814 578103 492842
rect 578069 492774 578103 492776
rect 578069 492742 578103 492774
rect 578069 492672 578103 492704
rect 578069 492670 578103 492672
rect 578069 492604 578103 492632
rect 578069 492598 578103 492604
rect 578069 492536 578103 492560
rect 578069 492526 578103 492536
rect 578069 492468 578103 492488
rect 578069 492454 578103 492468
rect 578069 492400 578103 492416
rect 578069 492382 578103 492400
rect 578069 492332 578103 492344
rect 578069 492310 578103 492332
rect 578069 492264 578103 492272
rect 578069 492238 578103 492264
rect 578327 493182 578361 493208
rect 578327 493174 578361 493182
rect 578327 493114 578361 493136
rect 578327 493102 578361 493114
rect 578327 493046 578361 493064
rect 578327 493030 578361 493046
rect 578327 492978 578361 492992
rect 578327 492958 578361 492978
rect 578327 492910 578361 492920
rect 578327 492886 578361 492910
rect 578327 492842 578361 492848
rect 578327 492814 578361 492842
rect 578327 492774 578361 492776
rect 578327 492742 578361 492774
rect 578327 492672 578361 492704
rect 578327 492670 578361 492672
rect 578327 492604 578361 492632
rect 578327 492598 578361 492604
rect 578327 492536 578361 492560
rect 578327 492526 578361 492536
rect 578327 492468 578361 492488
rect 578327 492454 578361 492468
rect 578327 492400 578361 492416
rect 578327 492382 578361 492400
rect 578327 492332 578361 492344
rect 578327 492310 578361 492332
rect 578327 492264 578361 492272
rect 578327 492238 578361 492264
rect 578585 493182 578619 493208
rect 578585 493174 578619 493182
rect 578585 493114 578619 493136
rect 578585 493102 578619 493114
rect 578585 493046 578619 493064
rect 578585 493030 578619 493046
rect 578585 492978 578619 492992
rect 578585 492958 578619 492978
rect 578585 492910 578619 492920
rect 578585 492886 578619 492910
rect 578585 492842 578619 492848
rect 578585 492814 578619 492842
rect 578585 492774 578619 492776
rect 578585 492742 578619 492774
rect 578585 492672 578619 492704
rect 578585 492670 578619 492672
rect 578585 492604 578619 492632
rect 578585 492598 578619 492604
rect 578585 492536 578619 492560
rect 578585 492526 578619 492536
rect 578585 492468 578619 492488
rect 578585 492454 578619 492468
rect 578585 492400 578619 492416
rect 578585 492382 578619 492400
rect 578585 492332 578619 492344
rect 578585 492310 578619 492332
rect 578585 492264 578619 492272
rect 578585 492238 578619 492264
rect 578843 493182 578877 493208
rect 578843 493174 578877 493182
rect 578843 493114 578877 493136
rect 578843 493102 578877 493114
rect 578843 493046 578877 493064
rect 578843 493030 578877 493046
rect 578843 492978 578877 492992
rect 578843 492958 578877 492978
rect 578843 492910 578877 492920
rect 578843 492886 578877 492910
rect 578843 492842 578877 492848
rect 578843 492814 578877 492842
rect 578843 492774 578877 492776
rect 578843 492742 578877 492774
rect 578843 492672 578877 492704
rect 578843 492670 578877 492672
rect 578843 492604 578877 492632
rect 578843 492598 578877 492604
rect 578843 492536 578877 492560
rect 578843 492526 578877 492536
rect 578843 492468 578877 492488
rect 578843 492454 578877 492468
rect 578843 492400 578877 492416
rect 578843 492382 578877 492400
rect 578843 492332 578877 492344
rect 578843 492310 578877 492332
rect 578843 492264 578877 492272
rect 578843 492238 578877 492264
rect 579101 493182 579135 493208
rect 579101 493174 579135 493182
rect 579101 493114 579135 493136
rect 579101 493102 579135 493114
rect 579101 493046 579135 493064
rect 579101 493030 579135 493046
rect 579101 492978 579135 492992
rect 579101 492958 579135 492978
rect 579101 492910 579135 492920
rect 579101 492886 579135 492910
rect 579101 492842 579135 492848
rect 579101 492814 579135 492842
rect 579101 492774 579135 492776
rect 579101 492742 579135 492774
rect 579101 492672 579135 492704
rect 579101 492670 579135 492672
rect 579101 492604 579135 492632
rect 579101 492598 579135 492604
rect 579101 492536 579135 492560
rect 579101 492526 579135 492536
rect 579101 492468 579135 492488
rect 579101 492454 579135 492468
rect 579101 492400 579135 492416
rect 579101 492382 579135 492400
rect 579101 492332 579135 492344
rect 579101 492310 579135 492332
rect 579101 492264 579135 492272
rect 579101 492238 579135 492264
rect 579359 493182 579393 493208
rect 579359 493174 579393 493182
rect 579359 493114 579393 493136
rect 579359 493102 579393 493114
rect 579359 493046 579393 493064
rect 579359 493030 579393 493046
rect 579359 492978 579393 492992
rect 579359 492958 579393 492978
rect 579359 492910 579393 492920
rect 579359 492886 579393 492910
rect 579359 492842 579393 492848
rect 579359 492814 579393 492842
rect 579359 492774 579393 492776
rect 579359 492742 579393 492774
rect 579359 492672 579393 492704
rect 579359 492670 579393 492672
rect 579359 492604 579393 492632
rect 579359 492598 579393 492604
rect 579359 492536 579393 492560
rect 579359 492526 579393 492536
rect 579359 492468 579393 492488
rect 579359 492454 579393 492468
rect 579359 492400 579393 492416
rect 579359 492382 579393 492400
rect 579359 492332 579393 492344
rect 579359 492310 579393 492332
rect 579359 492264 579393 492272
rect 579359 492238 579393 492264
rect 579617 493182 579651 493208
rect 579617 493174 579651 493182
rect 579617 493114 579651 493136
rect 579617 493102 579651 493114
rect 579617 493046 579651 493064
rect 579617 493030 579651 493046
rect 579617 492978 579651 492992
rect 579617 492958 579651 492978
rect 579617 492910 579651 492920
rect 579617 492886 579651 492910
rect 579617 492842 579651 492848
rect 579617 492814 579651 492842
rect 579617 492774 579651 492776
rect 579617 492742 579651 492774
rect 579617 492672 579651 492704
rect 579617 492670 579651 492672
rect 579617 492604 579651 492632
rect 579617 492598 579651 492604
rect 579617 492536 579651 492560
rect 579617 492526 579651 492536
rect 579617 492468 579651 492488
rect 579617 492454 579651 492468
rect 579617 492400 579651 492416
rect 579617 492382 579651 492400
rect 579617 492332 579651 492344
rect 579617 492310 579651 492332
rect 579617 492264 579651 492272
rect 579617 492238 579651 492264
rect 579875 493182 579909 493208
rect 579875 493174 579909 493182
rect 579875 493114 579909 493136
rect 579875 493102 579909 493114
rect 579875 493046 579909 493064
rect 579875 493030 579909 493046
rect 579875 492978 579909 492992
rect 579875 492958 579909 492978
rect 579875 492910 579909 492920
rect 579875 492886 579909 492910
rect 579875 492842 579909 492848
rect 579875 492814 579909 492842
rect 579875 492774 579909 492776
rect 579875 492742 579909 492774
rect 579875 492672 579909 492704
rect 579875 492670 579909 492672
rect 579875 492604 579909 492632
rect 579875 492598 579909 492604
rect 579875 492536 579909 492560
rect 579875 492526 579909 492536
rect 579875 492468 579909 492488
rect 579875 492454 579909 492468
rect 579875 492400 579909 492416
rect 579875 492382 579909 492400
rect 579875 492332 579909 492344
rect 579875 492310 579909 492332
rect 579875 492264 579909 492272
rect 579875 492238 579909 492264
rect 580133 493182 580167 493208
rect 580133 493174 580167 493182
rect 580133 493114 580167 493136
rect 580133 493102 580167 493114
rect 580133 493046 580167 493064
rect 580133 493030 580167 493046
rect 580133 492978 580167 492992
rect 580133 492958 580167 492978
rect 580133 492910 580167 492920
rect 580133 492886 580167 492910
rect 580133 492842 580167 492848
rect 580133 492814 580167 492842
rect 580133 492774 580167 492776
rect 580133 492742 580167 492774
rect 580133 492672 580167 492704
rect 580133 492670 580167 492672
rect 580133 492604 580167 492632
rect 580133 492598 580167 492604
rect 580133 492536 580167 492560
rect 580133 492526 580167 492536
rect 580133 492468 580167 492488
rect 580133 492454 580167 492468
rect 580133 492400 580167 492416
rect 580133 492382 580167 492400
rect 580133 492332 580167 492344
rect 580133 492310 580167 492332
rect 580133 492264 580167 492272
rect 580133 492238 580167 492264
rect 580391 493182 580425 493208
rect 580391 493174 580425 493182
rect 580391 493114 580425 493136
rect 580391 493102 580425 493114
rect 580391 493046 580425 493064
rect 580391 493030 580425 493046
rect 580391 492978 580425 492992
rect 580391 492958 580425 492978
rect 580391 492910 580425 492920
rect 580391 492886 580425 492910
rect 580391 492842 580425 492848
rect 580391 492814 580425 492842
rect 580391 492774 580425 492776
rect 580391 492742 580425 492774
rect 580391 492672 580425 492704
rect 580391 492670 580425 492672
rect 580391 492604 580425 492632
rect 580391 492598 580425 492604
rect 580391 492536 580425 492560
rect 580391 492526 580425 492536
rect 580391 492468 580425 492488
rect 580391 492454 580425 492468
rect 580391 492400 580425 492416
rect 580391 492382 580425 492400
rect 580391 492332 580425 492344
rect 580391 492310 580425 492332
rect 580391 492264 580425 492272
rect 580391 492238 580425 492264
rect 560863 491932 560897 491966
rect 561063 491932 561097 491966
rect 561263 491932 561297 491966
rect 561463 491932 561497 491966
rect 561663 491932 561697 491966
rect 561863 491932 561897 491966
rect 562063 491932 562097 491966
rect 562263 491932 562297 491966
rect 562463 491932 562497 491966
rect 562663 491932 562697 491966
rect 562863 491932 562897 491966
rect 563063 491932 563097 491966
rect 563263 491932 563297 491966
rect 563463 491932 563497 491966
rect 563663 491932 563697 491966
rect 563863 491932 563897 491966
rect 564063 491932 564097 491966
rect 564263 491932 564297 491966
rect 564463 491932 564497 491966
rect 564663 491932 564697 491966
rect 564863 491932 564897 491966
rect 565063 491932 565097 491966
rect 565263 491932 565297 491966
rect 565463 491932 565497 491966
rect 565663 491932 565697 491966
rect 580584 492066 580618 492100
rect 574977 491924 575011 491958
rect 575255 491706 575289 491740
rect 575455 491706 575489 491740
rect 575655 491706 575689 491740
rect 575855 491706 575889 491740
rect 576055 491706 576089 491740
rect 576255 491706 576289 491740
rect 576455 491706 576489 491740
rect 576655 491706 576689 491740
rect 576855 491706 576889 491740
rect 577055 491706 577089 491740
rect 577255 491706 577289 491740
rect 577455 491706 577489 491740
rect 577655 491706 577689 491740
rect 577855 491706 577889 491740
rect 578055 491706 578089 491740
rect 578255 491706 578289 491740
rect 578455 491706 578489 491740
rect 578655 491706 578689 491740
rect 578855 491706 578889 491740
rect 579055 491706 579089 491740
rect 579255 491706 579289 491740
rect 579455 491706 579489 491740
rect 579655 491706 579689 491740
rect 579855 491706 579889 491740
rect 580055 491706 580089 491740
rect 580255 491706 580289 491740
rect 560799 404670 560833 404704
rect 560999 404670 561033 404704
rect 561199 404670 561233 404704
rect 561399 404670 561433 404704
rect 561599 404670 561633 404704
rect 561799 404670 561833 404704
rect 561999 404670 562033 404704
rect 562199 404670 562233 404704
rect 562399 404670 562433 404704
rect 562599 404670 562633 404704
rect 562799 404670 562833 404704
rect 562999 404670 563033 404704
rect 563199 404670 563233 404704
rect 563399 404670 563433 404704
rect 563599 404670 563633 404704
rect 563799 404670 563833 404704
rect 563999 404670 564033 404704
rect 564199 404670 564233 404704
rect 564399 404670 564433 404704
rect 564599 404670 564633 404704
rect 564799 404670 564833 404704
rect 564999 404670 565033 404704
rect 565199 404670 565233 404704
rect 565399 404670 565433 404704
rect 565599 404670 565633 404704
rect 560303 403221 560409 403327
rect 560611 404266 560645 404292
rect 560611 404258 560645 404266
rect 560611 404198 560645 404220
rect 560611 404186 560645 404198
rect 560611 404130 560645 404148
rect 560611 404114 560645 404130
rect 560611 404062 560645 404076
rect 560611 404042 560645 404062
rect 560611 403994 560645 404004
rect 560611 403970 560645 403994
rect 560611 403926 560645 403932
rect 560611 403898 560645 403926
rect 560611 403858 560645 403860
rect 560611 403826 560645 403858
rect 560611 403756 560645 403788
rect 560611 403754 560645 403756
rect 560611 403688 560645 403716
rect 560611 403682 560645 403688
rect 560611 403620 560645 403644
rect 560611 403610 560645 403620
rect 560611 403552 560645 403572
rect 560611 403538 560645 403552
rect 560611 403484 560645 403500
rect 560611 403466 560645 403484
rect 560611 403416 560645 403428
rect 560611 403394 560645 403416
rect 560611 403348 560645 403356
rect 560611 403322 560645 403348
rect 560869 404266 560903 404292
rect 560869 404258 560903 404266
rect 560869 404198 560903 404220
rect 560869 404186 560903 404198
rect 560869 404130 560903 404148
rect 560869 404114 560903 404130
rect 560869 404062 560903 404076
rect 560869 404042 560903 404062
rect 560869 403994 560903 404004
rect 560869 403970 560903 403994
rect 560869 403926 560903 403932
rect 560869 403898 560903 403926
rect 560869 403858 560903 403860
rect 560869 403826 560903 403858
rect 560869 403756 560903 403788
rect 560869 403754 560903 403756
rect 560869 403688 560903 403716
rect 560869 403682 560903 403688
rect 560869 403620 560903 403644
rect 560869 403610 560903 403620
rect 560869 403552 560903 403572
rect 560869 403538 560903 403552
rect 560869 403484 560903 403500
rect 560869 403466 560903 403484
rect 560869 403416 560903 403428
rect 560869 403394 560903 403416
rect 560869 403348 560903 403356
rect 560869 403322 560903 403348
rect 561127 404266 561161 404292
rect 561127 404258 561161 404266
rect 561127 404198 561161 404220
rect 561127 404186 561161 404198
rect 561127 404130 561161 404148
rect 561127 404114 561161 404130
rect 561127 404062 561161 404076
rect 561127 404042 561161 404062
rect 561127 403994 561161 404004
rect 561127 403970 561161 403994
rect 561127 403926 561161 403932
rect 561127 403898 561161 403926
rect 561127 403858 561161 403860
rect 561127 403826 561161 403858
rect 561127 403756 561161 403788
rect 561127 403754 561161 403756
rect 561127 403688 561161 403716
rect 561127 403682 561161 403688
rect 561127 403620 561161 403644
rect 561127 403610 561161 403620
rect 561127 403552 561161 403572
rect 561127 403538 561161 403552
rect 561127 403484 561161 403500
rect 561127 403466 561161 403484
rect 561127 403416 561161 403428
rect 561127 403394 561161 403416
rect 561127 403348 561161 403356
rect 561127 403322 561161 403348
rect 561385 404266 561419 404292
rect 561385 404258 561419 404266
rect 561385 404198 561419 404220
rect 561385 404186 561419 404198
rect 561385 404130 561419 404148
rect 561385 404114 561419 404130
rect 561385 404062 561419 404076
rect 561385 404042 561419 404062
rect 561385 403994 561419 404004
rect 561385 403970 561419 403994
rect 561385 403926 561419 403932
rect 561385 403898 561419 403926
rect 561385 403858 561419 403860
rect 561385 403826 561419 403858
rect 561385 403756 561419 403788
rect 561385 403754 561419 403756
rect 561385 403688 561419 403716
rect 561385 403682 561419 403688
rect 561385 403620 561419 403644
rect 561385 403610 561419 403620
rect 561385 403552 561419 403572
rect 561385 403538 561419 403552
rect 561385 403484 561419 403500
rect 561385 403466 561419 403484
rect 561385 403416 561419 403428
rect 561385 403394 561419 403416
rect 561385 403348 561419 403356
rect 561385 403322 561419 403348
rect 561643 404266 561677 404292
rect 561643 404258 561677 404266
rect 561643 404198 561677 404220
rect 561643 404186 561677 404198
rect 561643 404130 561677 404148
rect 561643 404114 561677 404130
rect 561643 404062 561677 404076
rect 561643 404042 561677 404062
rect 561643 403994 561677 404004
rect 561643 403970 561677 403994
rect 561643 403926 561677 403932
rect 561643 403898 561677 403926
rect 561643 403858 561677 403860
rect 561643 403826 561677 403858
rect 561643 403756 561677 403788
rect 561643 403754 561677 403756
rect 561643 403688 561677 403716
rect 561643 403682 561677 403688
rect 561643 403620 561677 403644
rect 561643 403610 561677 403620
rect 561643 403552 561677 403572
rect 561643 403538 561677 403552
rect 561643 403484 561677 403500
rect 561643 403466 561677 403484
rect 561643 403416 561677 403428
rect 561643 403394 561677 403416
rect 561643 403348 561677 403356
rect 561643 403322 561677 403348
rect 561901 404266 561935 404292
rect 561901 404258 561935 404266
rect 561901 404198 561935 404220
rect 561901 404186 561935 404198
rect 561901 404130 561935 404148
rect 561901 404114 561935 404130
rect 561901 404062 561935 404076
rect 561901 404042 561935 404062
rect 561901 403994 561935 404004
rect 561901 403970 561935 403994
rect 561901 403926 561935 403932
rect 561901 403898 561935 403926
rect 561901 403858 561935 403860
rect 561901 403826 561935 403858
rect 561901 403756 561935 403788
rect 561901 403754 561935 403756
rect 561901 403688 561935 403716
rect 561901 403682 561935 403688
rect 561901 403620 561935 403644
rect 561901 403610 561935 403620
rect 561901 403552 561935 403572
rect 561901 403538 561935 403552
rect 561901 403484 561935 403500
rect 561901 403466 561935 403484
rect 561901 403416 561935 403428
rect 561901 403394 561935 403416
rect 561901 403348 561935 403356
rect 561901 403322 561935 403348
rect 562159 404266 562193 404292
rect 562159 404258 562193 404266
rect 562159 404198 562193 404220
rect 562159 404186 562193 404198
rect 562159 404130 562193 404148
rect 562159 404114 562193 404130
rect 562159 404062 562193 404076
rect 562159 404042 562193 404062
rect 562159 403994 562193 404004
rect 562159 403970 562193 403994
rect 562159 403926 562193 403932
rect 562159 403898 562193 403926
rect 562159 403858 562193 403860
rect 562159 403826 562193 403858
rect 562159 403756 562193 403788
rect 562159 403754 562193 403756
rect 562159 403688 562193 403716
rect 562159 403682 562193 403688
rect 562159 403620 562193 403644
rect 562159 403610 562193 403620
rect 562159 403552 562193 403572
rect 562159 403538 562193 403552
rect 562159 403484 562193 403500
rect 562159 403466 562193 403484
rect 562159 403416 562193 403428
rect 562159 403394 562193 403416
rect 562159 403348 562193 403356
rect 562159 403322 562193 403348
rect 562417 404266 562451 404292
rect 562417 404258 562451 404266
rect 562417 404198 562451 404220
rect 562417 404186 562451 404198
rect 562417 404130 562451 404148
rect 562417 404114 562451 404130
rect 562417 404062 562451 404076
rect 562417 404042 562451 404062
rect 562417 403994 562451 404004
rect 562417 403970 562451 403994
rect 562417 403926 562451 403932
rect 562417 403898 562451 403926
rect 562417 403858 562451 403860
rect 562417 403826 562451 403858
rect 562417 403756 562451 403788
rect 562417 403754 562451 403756
rect 562417 403688 562451 403716
rect 562417 403682 562451 403688
rect 562417 403620 562451 403644
rect 562417 403610 562451 403620
rect 562417 403552 562451 403572
rect 562417 403538 562451 403552
rect 562417 403484 562451 403500
rect 562417 403466 562451 403484
rect 562417 403416 562451 403428
rect 562417 403394 562451 403416
rect 562417 403348 562451 403356
rect 562417 403322 562451 403348
rect 562675 404266 562709 404292
rect 562675 404258 562709 404266
rect 562675 404198 562709 404220
rect 562675 404186 562709 404198
rect 562675 404130 562709 404148
rect 562675 404114 562709 404130
rect 562675 404062 562709 404076
rect 562675 404042 562709 404062
rect 562675 403994 562709 404004
rect 562675 403970 562709 403994
rect 562675 403926 562709 403932
rect 562675 403898 562709 403926
rect 562675 403858 562709 403860
rect 562675 403826 562709 403858
rect 562675 403756 562709 403788
rect 562675 403754 562709 403756
rect 562675 403688 562709 403716
rect 562675 403682 562709 403688
rect 562675 403620 562709 403644
rect 562675 403610 562709 403620
rect 562675 403552 562709 403572
rect 562675 403538 562709 403552
rect 562675 403484 562709 403500
rect 562675 403466 562709 403484
rect 562675 403416 562709 403428
rect 562675 403394 562709 403416
rect 562675 403348 562709 403356
rect 562675 403322 562709 403348
rect 562933 404266 562967 404292
rect 562933 404258 562967 404266
rect 562933 404198 562967 404220
rect 562933 404186 562967 404198
rect 562933 404130 562967 404148
rect 562933 404114 562967 404130
rect 562933 404062 562967 404076
rect 562933 404042 562967 404062
rect 562933 403994 562967 404004
rect 562933 403970 562967 403994
rect 562933 403926 562967 403932
rect 562933 403898 562967 403926
rect 562933 403858 562967 403860
rect 562933 403826 562967 403858
rect 562933 403756 562967 403788
rect 562933 403754 562967 403756
rect 562933 403688 562967 403716
rect 562933 403682 562967 403688
rect 562933 403620 562967 403644
rect 562933 403610 562967 403620
rect 562933 403552 562967 403572
rect 562933 403538 562967 403552
rect 562933 403484 562967 403500
rect 562933 403466 562967 403484
rect 562933 403416 562967 403428
rect 562933 403394 562967 403416
rect 562933 403348 562967 403356
rect 562933 403322 562967 403348
rect 563191 404266 563225 404292
rect 563191 404258 563225 404266
rect 563191 404198 563225 404220
rect 563191 404186 563225 404198
rect 563191 404130 563225 404148
rect 563191 404114 563225 404130
rect 563191 404062 563225 404076
rect 563191 404042 563225 404062
rect 563191 403994 563225 404004
rect 563191 403970 563225 403994
rect 563191 403926 563225 403932
rect 563191 403898 563225 403926
rect 563191 403858 563225 403860
rect 563191 403826 563225 403858
rect 563191 403756 563225 403788
rect 563191 403754 563225 403756
rect 563191 403688 563225 403716
rect 563191 403682 563225 403688
rect 563191 403620 563225 403644
rect 563191 403610 563225 403620
rect 563191 403552 563225 403572
rect 563191 403538 563225 403552
rect 563191 403484 563225 403500
rect 563191 403466 563225 403484
rect 563191 403416 563225 403428
rect 563191 403394 563225 403416
rect 563191 403348 563225 403356
rect 563191 403322 563225 403348
rect 563449 404266 563483 404292
rect 563449 404258 563483 404266
rect 563449 404198 563483 404220
rect 563449 404186 563483 404198
rect 563449 404130 563483 404148
rect 563449 404114 563483 404130
rect 563449 404062 563483 404076
rect 563449 404042 563483 404062
rect 563449 403994 563483 404004
rect 563449 403970 563483 403994
rect 563449 403926 563483 403932
rect 563449 403898 563483 403926
rect 563449 403858 563483 403860
rect 563449 403826 563483 403858
rect 563449 403756 563483 403788
rect 563449 403754 563483 403756
rect 563449 403688 563483 403716
rect 563449 403682 563483 403688
rect 563449 403620 563483 403644
rect 563449 403610 563483 403620
rect 563449 403552 563483 403572
rect 563449 403538 563483 403552
rect 563449 403484 563483 403500
rect 563449 403466 563483 403484
rect 563449 403416 563483 403428
rect 563449 403394 563483 403416
rect 563449 403348 563483 403356
rect 563449 403322 563483 403348
rect 563707 404266 563741 404292
rect 563707 404258 563741 404266
rect 563707 404198 563741 404220
rect 563707 404186 563741 404198
rect 563707 404130 563741 404148
rect 563707 404114 563741 404130
rect 563707 404062 563741 404076
rect 563707 404042 563741 404062
rect 563707 403994 563741 404004
rect 563707 403970 563741 403994
rect 563707 403926 563741 403932
rect 563707 403898 563741 403926
rect 563707 403858 563741 403860
rect 563707 403826 563741 403858
rect 563707 403756 563741 403788
rect 563707 403754 563741 403756
rect 563707 403688 563741 403716
rect 563707 403682 563741 403688
rect 563707 403620 563741 403644
rect 563707 403610 563741 403620
rect 563707 403552 563741 403572
rect 563707 403538 563741 403552
rect 563707 403484 563741 403500
rect 563707 403466 563741 403484
rect 563707 403416 563741 403428
rect 563707 403394 563741 403416
rect 563707 403348 563741 403356
rect 563707 403322 563741 403348
rect 563965 404266 563999 404292
rect 563965 404258 563999 404266
rect 563965 404198 563999 404220
rect 563965 404186 563999 404198
rect 563965 404130 563999 404148
rect 563965 404114 563999 404130
rect 563965 404062 563999 404076
rect 563965 404042 563999 404062
rect 563965 403994 563999 404004
rect 563965 403970 563999 403994
rect 563965 403926 563999 403932
rect 563965 403898 563999 403926
rect 563965 403858 563999 403860
rect 563965 403826 563999 403858
rect 563965 403756 563999 403788
rect 563965 403754 563999 403756
rect 563965 403688 563999 403716
rect 563965 403682 563999 403688
rect 563965 403620 563999 403644
rect 563965 403610 563999 403620
rect 563965 403552 563999 403572
rect 563965 403538 563999 403552
rect 563965 403484 563999 403500
rect 563965 403466 563999 403484
rect 563965 403416 563999 403428
rect 563965 403394 563999 403416
rect 563965 403348 563999 403356
rect 563965 403322 563999 403348
rect 564223 404266 564257 404292
rect 564223 404258 564257 404266
rect 564223 404198 564257 404220
rect 564223 404186 564257 404198
rect 564223 404130 564257 404148
rect 564223 404114 564257 404130
rect 564223 404062 564257 404076
rect 564223 404042 564257 404062
rect 564223 403994 564257 404004
rect 564223 403970 564257 403994
rect 564223 403926 564257 403932
rect 564223 403898 564257 403926
rect 564223 403858 564257 403860
rect 564223 403826 564257 403858
rect 564223 403756 564257 403788
rect 564223 403754 564257 403756
rect 564223 403688 564257 403716
rect 564223 403682 564257 403688
rect 564223 403620 564257 403644
rect 564223 403610 564257 403620
rect 564223 403552 564257 403572
rect 564223 403538 564257 403552
rect 564223 403484 564257 403500
rect 564223 403466 564257 403484
rect 564223 403416 564257 403428
rect 564223 403394 564257 403416
rect 564223 403348 564257 403356
rect 564223 403322 564257 403348
rect 564481 404266 564515 404292
rect 564481 404258 564515 404266
rect 564481 404198 564515 404220
rect 564481 404186 564515 404198
rect 564481 404130 564515 404148
rect 564481 404114 564515 404130
rect 564481 404062 564515 404076
rect 564481 404042 564515 404062
rect 564481 403994 564515 404004
rect 564481 403970 564515 403994
rect 564481 403926 564515 403932
rect 564481 403898 564515 403926
rect 564481 403858 564515 403860
rect 564481 403826 564515 403858
rect 564481 403756 564515 403788
rect 564481 403754 564515 403756
rect 564481 403688 564515 403716
rect 564481 403682 564515 403688
rect 564481 403620 564515 403644
rect 564481 403610 564515 403620
rect 564481 403552 564515 403572
rect 564481 403538 564515 403552
rect 564481 403484 564515 403500
rect 564481 403466 564515 403484
rect 564481 403416 564515 403428
rect 564481 403394 564515 403416
rect 564481 403348 564515 403356
rect 564481 403322 564515 403348
rect 564739 404266 564773 404292
rect 564739 404258 564773 404266
rect 564739 404198 564773 404220
rect 564739 404186 564773 404198
rect 564739 404130 564773 404148
rect 564739 404114 564773 404130
rect 564739 404062 564773 404076
rect 564739 404042 564773 404062
rect 564739 403994 564773 404004
rect 564739 403970 564773 403994
rect 564739 403926 564773 403932
rect 564739 403898 564773 403926
rect 564739 403858 564773 403860
rect 564739 403826 564773 403858
rect 564739 403756 564773 403788
rect 564739 403754 564773 403756
rect 564739 403688 564773 403716
rect 564739 403682 564773 403688
rect 564739 403620 564773 403644
rect 564739 403610 564773 403620
rect 564739 403552 564773 403572
rect 564739 403538 564773 403552
rect 564739 403484 564773 403500
rect 564739 403466 564773 403484
rect 564739 403416 564773 403428
rect 564739 403394 564773 403416
rect 564739 403348 564773 403356
rect 564739 403322 564773 403348
rect 564997 404266 565031 404292
rect 564997 404258 565031 404266
rect 564997 404198 565031 404220
rect 564997 404186 565031 404198
rect 564997 404130 565031 404148
rect 564997 404114 565031 404130
rect 564997 404062 565031 404076
rect 564997 404042 565031 404062
rect 564997 403994 565031 404004
rect 564997 403970 565031 403994
rect 564997 403926 565031 403932
rect 564997 403898 565031 403926
rect 564997 403858 565031 403860
rect 564997 403826 565031 403858
rect 564997 403756 565031 403788
rect 564997 403754 565031 403756
rect 564997 403688 565031 403716
rect 564997 403682 565031 403688
rect 564997 403620 565031 403644
rect 564997 403610 565031 403620
rect 564997 403552 565031 403572
rect 564997 403538 565031 403552
rect 564997 403484 565031 403500
rect 564997 403466 565031 403484
rect 564997 403416 565031 403428
rect 564997 403394 565031 403416
rect 564997 403348 565031 403356
rect 564997 403322 565031 403348
rect 565255 404266 565289 404292
rect 565255 404258 565289 404266
rect 565255 404198 565289 404220
rect 565255 404186 565289 404198
rect 565255 404130 565289 404148
rect 565255 404114 565289 404130
rect 565255 404062 565289 404076
rect 565255 404042 565289 404062
rect 565255 403994 565289 404004
rect 565255 403970 565289 403994
rect 565255 403926 565289 403932
rect 565255 403898 565289 403926
rect 565255 403858 565289 403860
rect 565255 403826 565289 403858
rect 565255 403756 565289 403788
rect 565255 403754 565289 403756
rect 565255 403688 565289 403716
rect 565255 403682 565289 403688
rect 565255 403620 565289 403644
rect 565255 403610 565289 403620
rect 565255 403552 565289 403572
rect 565255 403538 565289 403552
rect 565255 403484 565289 403500
rect 565255 403466 565289 403484
rect 565255 403416 565289 403428
rect 565255 403394 565289 403416
rect 565255 403348 565289 403356
rect 565255 403322 565289 403348
rect 565513 404266 565547 404292
rect 565513 404258 565547 404266
rect 565513 404198 565547 404220
rect 565513 404186 565547 404198
rect 565513 404130 565547 404148
rect 565513 404114 565547 404130
rect 565513 404062 565547 404076
rect 565513 404042 565547 404062
rect 565513 403994 565547 404004
rect 565513 403970 565547 403994
rect 565513 403926 565547 403932
rect 565513 403898 565547 403926
rect 565513 403858 565547 403860
rect 565513 403826 565547 403858
rect 565513 403756 565547 403788
rect 565513 403754 565547 403756
rect 565513 403688 565547 403716
rect 565513 403682 565547 403688
rect 565513 403620 565547 403644
rect 565513 403610 565547 403620
rect 565513 403552 565547 403572
rect 565513 403538 565547 403552
rect 565513 403484 565547 403500
rect 565513 403466 565547 403484
rect 565513 403416 565547 403428
rect 565513 403394 565547 403416
rect 565513 403348 565547 403356
rect 565513 403322 565547 403348
rect 565771 404266 565805 404292
rect 565771 404258 565805 404266
rect 565771 404198 565805 404220
rect 565771 404186 565805 404198
rect 565771 404130 565805 404148
rect 565771 404114 565805 404130
rect 565771 404062 565805 404076
rect 565771 404042 565805 404062
rect 565771 403994 565805 404004
rect 565771 403970 565805 403994
rect 565771 403926 565805 403932
rect 565771 403898 565805 403926
rect 565771 403858 565805 403860
rect 565771 403826 565805 403858
rect 565771 403756 565805 403788
rect 565771 403754 565805 403756
rect 565771 403688 565805 403716
rect 565771 403682 565805 403688
rect 565771 403620 565805 403644
rect 565771 403610 565805 403620
rect 565771 403552 565805 403572
rect 565771 403538 565805 403552
rect 565771 403484 565805 403500
rect 565771 403466 565805 403484
rect 565771 403416 565805 403428
rect 565771 403394 565805 403416
rect 565771 403348 565805 403356
rect 565771 403322 565805 403348
rect 566051 403188 566157 403294
rect 560799 402790 560833 402824
rect 560999 402790 561033 402824
rect 561199 402790 561233 402824
rect 561399 402790 561433 402824
rect 561599 402790 561633 402824
rect 561799 402790 561833 402824
rect 561999 402790 562033 402824
rect 562199 402790 562233 402824
rect 562399 402790 562433 402824
rect 562599 402790 562633 402824
rect 562799 402790 562833 402824
rect 562999 402790 563033 402824
rect 563199 402790 563233 402824
rect 563399 402790 563433 402824
rect 563599 402790 563633 402824
rect 563799 402790 563833 402824
rect 563999 402790 564033 402824
rect 564199 402790 564233 402824
rect 564399 402790 564433 402824
rect 564599 402790 564633 402824
rect 564799 402790 564833 402824
rect 564999 402790 565033 402824
rect 565199 402790 565233 402824
rect 565399 402790 565433 402824
rect 565599 402790 565633 402824
rect 560755 359352 560789 359386
rect 560955 359352 560989 359386
rect 561155 359352 561189 359386
rect 561355 359352 561389 359386
rect 561555 359352 561589 359386
rect 561755 359352 561789 359386
rect 561955 359352 561989 359386
rect 562155 359352 562189 359386
rect 562355 359352 562389 359386
rect 562555 359352 562589 359386
rect 562755 359352 562789 359386
rect 562955 359352 562989 359386
rect 563155 359352 563189 359386
rect 563355 359352 563389 359386
rect 563555 359352 563589 359386
rect 563755 359352 563789 359386
rect 563955 359352 563989 359386
rect 564155 359352 564189 359386
rect 564355 359352 564389 359386
rect 564555 359352 564589 359386
rect 564755 359352 564789 359386
rect 564955 359352 564989 359386
rect 565155 359352 565189 359386
rect 565355 359352 565389 359386
rect 565555 359352 565589 359386
rect 574729 359282 574763 359316
rect 574929 359282 574963 359316
rect 575129 359282 575163 359316
rect 575329 359282 575363 359316
rect 575529 359282 575563 359316
rect 575729 359282 575763 359316
rect 575929 359282 575963 359316
rect 576129 359282 576163 359316
rect 576329 359282 576363 359316
rect 576529 359282 576563 359316
rect 576729 359282 576763 359316
rect 576929 359282 576963 359316
rect 577129 359282 577163 359316
rect 577329 359282 577363 359316
rect 577529 359282 577563 359316
rect 577729 359282 577763 359316
rect 577929 359282 577963 359316
rect 578129 359282 578163 359316
rect 578329 359282 578363 359316
rect 578529 359282 578563 359316
rect 578729 359282 578763 359316
rect 578929 359282 578963 359316
rect 579129 359282 579163 359316
rect 579329 359282 579363 359316
rect 579529 359282 579563 359316
rect 579729 359282 579763 359316
rect 560259 357903 560365 358009
rect 560567 358948 560601 358974
rect 560567 358940 560601 358948
rect 560567 358880 560601 358902
rect 560567 358868 560601 358880
rect 560567 358812 560601 358830
rect 560567 358796 560601 358812
rect 560567 358744 560601 358758
rect 560567 358724 560601 358744
rect 560567 358676 560601 358686
rect 560567 358652 560601 358676
rect 560567 358608 560601 358614
rect 560567 358580 560601 358608
rect 560567 358540 560601 358542
rect 560567 358508 560601 358540
rect 560567 358438 560601 358470
rect 560567 358436 560601 358438
rect 560567 358370 560601 358398
rect 560567 358364 560601 358370
rect 560567 358302 560601 358326
rect 560567 358292 560601 358302
rect 560567 358234 560601 358254
rect 560567 358220 560601 358234
rect 560567 358166 560601 358182
rect 560567 358148 560601 358166
rect 560567 358098 560601 358110
rect 560567 358076 560601 358098
rect 560567 358030 560601 358038
rect 560567 358004 560601 358030
rect 560825 358948 560859 358974
rect 560825 358940 560859 358948
rect 560825 358880 560859 358902
rect 560825 358868 560859 358880
rect 560825 358812 560859 358830
rect 560825 358796 560859 358812
rect 560825 358744 560859 358758
rect 560825 358724 560859 358744
rect 560825 358676 560859 358686
rect 560825 358652 560859 358676
rect 560825 358608 560859 358614
rect 560825 358580 560859 358608
rect 560825 358540 560859 358542
rect 560825 358508 560859 358540
rect 560825 358438 560859 358470
rect 560825 358436 560859 358438
rect 560825 358370 560859 358398
rect 560825 358364 560859 358370
rect 560825 358302 560859 358326
rect 560825 358292 560859 358302
rect 560825 358234 560859 358254
rect 560825 358220 560859 358234
rect 560825 358166 560859 358182
rect 560825 358148 560859 358166
rect 560825 358098 560859 358110
rect 560825 358076 560859 358098
rect 560825 358030 560859 358038
rect 560825 358004 560859 358030
rect 561083 358948 561117 358974
rect 561083 358940 561117 358948
rect 561083 358880 561117 358902
rect 561083 358868 561117 358880
rect 561083 358812 561117 358830
rect 561083 358796 561117 358812
rect 561083 358744 561117 358758
rect 561083 358724 561117 358744
rect 561083 358676 561117 358686
rect 561083 358652 561117 358676
rect 561083 358608 561117 358614
rect 561083 358580 561117 358608
rect 561083 358540 561117 358542
rect 561083 358508 561117 358540
rect 561083 358438 561117 358470
rect 561083 358436 561117 358438
rect 561083 358370 561117 358398
rect 561083 358364 561117 358370
rect 561083 358302 561117 358326
rect 561083 358292 561117 358302
rect 561083 358234 561117 358254
rect 561083 358220 561117 358234
rect 561083 358166 561117 358182
rect 561083 358148 561117 358166
rect 561083 358098 561117 358110
rect 561083 358076 561117 358098
rect 561083 358030 561117 358038
rect 561083 358004 561117 358030
rect 561341 358948 561375 358974
rect 561341 358940 561375 358948
rect 561341 358880 561375 358902
rect 561341 358868 561375 358880
rect 561341 358812 561375 358830
rect 561341 358796 561375 358812
rect 561341 358744 561375 358758
rect 561341 358724 561375 358744
rect 561341 358676 561375 358686
rect 561341 358652 561375 358676
rect 561341 358608 561375 358614
rect 561341 358580 561375 358608
rect 561341 358540 561375 358542
rect 561341 358508 561375 358540
rect 561341 358438 561375 358470
rect 561341 358436 561375 358438
rect 561341 358370 561375 358398
rect 561341 358364 561375 358370
rect 561341 358302 561375 358326
rect 561341 358292 561375 358302
rect 561341 358234 561375 358254
rect 561341 358220 561375 358234
rect 561341 358166 561375 358182
rect 561341 358148 561375 358166
rect 561341 358098 561375 358110
rect 561341 358076 561375 358098
rect 561341 358030 561375 358038
rect 561341 358004 561375 358030
rect 561599 358948 561633 358974
rect 561599 358940 561633 358948
rect 561599 358880 561633 358902
rect 561599 358868 561633 358880
rect 561599 358812 561633 358830
rect 561599 358796 561633 358812
rect 561599 358744 561633 358758
rect 561599 358724 561633 358744
rect 561599 358676 561633 358686
rect 561599 358652 561633 358676
rect 561599 358608 561633 358614
rect 561599 358580 561633 358608
rect 561599 358540 561633 358542
rect 561599 358508 561633 358540
rect 561599 358438 561633 358470
rect 561599 358436 561633 358438
rect 561599 358370 561633 358398
rect 561599 358364 561633 358370
rect 561599 358302 561633 358326
rect 561599 358292 561633 358302
rect 561599 358234 561633 358254
rect 561599 358220 561633 358234
rect 561599 358166 561633 358182
rect 561599 358148 561633 358166
rect 561599 358098 561633 358110
rect 561599 358076 561633 358098
rect 561599 358030 561633 358038
rect 561599 358004 561633 358030
rect 561857 358948 561891 358974
rect 561857 358940 561891 358948
rect 561857 358880 561891 358902
rect 561857 358868 561891 358880
rect 561857 358812 561891 358830
rect 561857 358796 561891 358812
rect 561857 358744 561891 358758
rect 561857 358724 561891 358744
rect 561857 358676 561891 358686
rect 561857 358652 561891 358676
rect 561857 358608 561891 358614
rect 561857 358580 561891 358608
rect 561857 358540 561891 358542
rect 561857 358508 561891 358540
rect 561857 358438 561891 358470
rect 561857 358436 561891 358438
rect 561857 358370 561891 358398
rect 561857 358364 561891 358370
rect 561857 358302 561891 358326
rect 561857 358292 561891 358302
rect 561857 358234 561891 358254
rect 561857 358220 561891 358234
rect 561857 358166 561891 358182
rect 561857 358148 561891 358166
rect 561857 358098 561891 358110
rect 561857 358076 561891 358098
rect 561857 358030 561891 358038
rect 561857 358004 561891 358030
rect 562115 358948 562149 358974
rect 562115 358940 562149 358948
rect 562115 358880 562149 358902
rect 562115 358868 562149 358880
rect 562115 358812 562149 358830
rect 562115 358796 562149 358812
rect 562115 358744 562149 358758
rect 562115 358724 562149 358744
rect 562115 358676 562149 358686
rect 562115 358652 562149 358676
rect 562115 358608 562149 358614
rect 562115 358580 562149 358608
rect 562115 358540 562149 358542
rect 562115 358508 562149 358540
rect 562115 358438 562149 358470
rect 562115 358436 562149 358438
rect 562115 358370 562149 358398
rect 562115 358364 562149 358370
rect 562115 358302 562149 358326
rect 562115 358292 562149 358302
rect 562115 358234 562149 358254
rect 562115 358220 562149 358234
rect 562115 358166 562149 358182
rect 562115 358148 562149 358166
rect 562115 358098 562149 358110
rect 562115 358076 562149 358098
rect 562115 358030 562149 358038
rect 562115 358004 562149 358030
rect 562373 358948 562407 358974
rect 562373 358940 562407 358948
rect 562373 358880 562407 358902
rect 562373 358868 562407 358880
rect 562373 358812 562407 358830
rect 562373 358796 562407 358812
rect 562373 358744 562407 358758
rect 562373 358724 562407 358744
rect 562373 358676 562407 358686
rect 562373 358652 562407 358676
rect 562373 358608 562407 358614
rect 562373 358580 562407 358608
rect 562373 358540 562407 358542
rect 562373 358508 562407 358540
rect 562373 358438 562407 358470
rect 562373 358436 562407 358438
rect 562373 358370 562407 358398
rect 562373 358364 562407 358370
rect 562373 358302 562407 358326
rect 562373 358292 562407 358302
rect 562373 358234 562407 358254
rect 562373 358220 562407 358234
rect 562373 358166 562407 358182
rect 562373 358148 562407 358166
rect 562373 358098 562407 358110
rect 562373 358076 562407 358098
rect 562373 358030 562407 358038
rect 562373 358004 562407 358030
rect 562631 358948 562665 358974
rect 562631 358940 562665 358948
rect 562631 358880 562665 358902
rect 562631 358868 562665 358880
rect 562631 358812 562665 358830
rect 562631 358796 562665 358812
rect 562631 358744 562665 358758
rect 562631 358724 562665 358744
rect 562631 358676 562665 358686
rect 562631 358652 562665 358676
rect 562631 358608 562665 358614
rect 562631 358580 562665 358608
rect 562631 358540 562665 358542
rect 562631 358508 562665 358540
rect 562631 358438 562665 358470
rect 562631 358436 562665 358438
rect 562631 358370 562665 358398
rect 562631 358364 562665 358370
rect 562631 358302 562665 358326
rect 562631 358292 562665 358302
rect 562631 358234 562665 358254
rect 562631 358220 562665 358234
rect 562631 358166 562665 358182
rect 562631 358148 562665 358166
rect 562631 358098 562665 358110
rect 562631 358076 562665 358098
rect 562631 358030 562665 358038
rect 562631 358004 562665 358030
rect 562889 358948 562923 358974
rect 562889 358940 562923 358948
rect 562889 358880 562923 358902
rect 562889 358868 562923 358880
rect 562889 358812 562923 358830
rect 562889 358796 562923 358812
rect 562889 358744 562923 358758
rect 562889 358724 562923 358744
rect 562889 358676 562923 358686
rect 562889 358652 562923 358676
rect 562889 358608 562923 358614
rect 562889 358580 562923 358608
rect 562889 358540 562923 358542
rect 562889 358508 562923 358540
rect 562889 358438 562923 358470
rect 562889 358436 562923 358438
rect 562889 358370 562923 358398
rect 562889 358364 562923 358370
rect 562889 358302 562923 358326
rect 562889 358292 562923 358302
rect 562889 358234 562923 358254
rect 562889 358220 562923 358234
rect 562889 358166 562923 358182
rect 562889 358148 562923 358166
rect 562889 358098 562923 358110
rect 562889 358076 562923 358098
rect 562889 358030 562923 358038
rect 562889 358004 562923 358030
rect 563147 358948 563181 358974
rect 563147 358940 563181 358948
rect 563147 358880 563181 358902
rect 563147 358868 563181 358880
rect 563147 358812 563181 358830
rect 563147 358796 563181 358812
rect 563147 358744 563181 358758
rect 563147 358724 563181 358744
rect 563147 358676 563181 358686
rect 563147 358652 563181 358676
rect 563147 358608 563181 358614
rect 563147 358580 563181 358608
rect 563147 358540 563181 358542
rect 563147 358508 563181 358540
rect 563147 358438 563181 358470
rect 563147 358436 563181 358438
rect 563147 358370 563181 358398
rect 563147 358364 563181 358370
rect 563147 358302 563181 358326
rect 563147 358292 563181 358302
rect 563147 358234 563181 358254
rect 563147 358220 563181 358234
rect 563147 358166 563181 358182
rect 563147 358148 563181 358166
rect 563147 358098 563181 358110
rect 563147 358076 563181 358098
rect 563147 358030 563181 358038
rect 563147 358004 563181 358030
rect 563405 358948 563439 358974
rect 563405 358940 563439 358948
rect 563405 358880 563439 358902
rect 563405 358868 563439 358880
rect 563405 358812 563439 358830
rect 563405 358796 563439 358812
rect 563405 358744 563439 358758
rect 563405 358724 563439 358744
rect 563405 358676 563439 358686
rect 563405 358652 563439 358676
rect 563405 358608 563439 358614
rect 563405 358580 563439 358608
rect 563405 358540 563439 358542
rect 563405 358508 563439 358540
rect 563405 358438 563439 358470
rect 563405 358436 563439 358438
rect 563405 358370 563439 358398
rect 563405 358364 563439 358370
rect 563405 358302 563439 358326
rect 563405 358292 563439 358302
rect 563405 358234 563439 358254
rect 563405 358220 563439 358234
rect 563405 358166 563439 358182
rect 563405 358148 563439 358166
rect 563405 358098 563439 358110
rect 563405 358076 563439 358098
rect 563405 358030 563439 358038
rect 563405 358004 563439 358030
rect 563663 358948 563697 358974
rect 563663 358940 563697 358948
rect 563663 358880 563697 358902
rect 563663 358868 563697 358880
rect 563663 358812 563697 358830
rect 563663 358796 563697 358812
rect 563663 358744 563697 358758
rect 563663 358724 563697 358744
rect 563663 358676 563697 358686
rect 563663 358652 563697 358676
rect 563663 358608 563697 358614
rect 563663 358580 563697 358608
rect 563663 358540 563697 358542
rect 563663 358508 563697 358540
rect 563663 358438 563697 358470
rect 563663 358436 563697 358438
rect 563663 358370 563697 358398
rect 563663 358364 563697 358370
rect 563663 358302 563697 358326
rect 563663 358292 563697 358302
rect 563663 358234 563697 358254
rect 563663 358220 563697 358234
rect 563663 358166 563697 358182
rect 563663 358148 563697 358166
rect 563663 358098 563697 358110
rect 563663 358076 563697 358098
rect 563663 358030 563697 358038
rect 563663 358004 563697 358030
rect 563921 358948 563955 358974
rect 563921 358940 563955 358948
rect 563921 358880 563955 358902
rect 563921 358868 563955 358880
rect 563921 358812 563955 358830
rect 563921 358796 563955 358812
rect 563921 358744 563955 358758
rect 563921 358724 563955 358744
rect 563921 358676 563955 358686
rect 563921 358652 563955 358676
rect 563921 358608 563955 358614
rect 563921 358580 563955 358608
rect 563921 358540 563955 358542
rect 563921 358508 563955 358540
rect 563921 358438 563955 358470
rect 563921 358436 563955 358438
rect 563921 358370 563955 358398
rect 563921 358364 563955 358370
rect 563921 358302 563955 358326
rect 563921 358292 563955 358302
rect 563921 358234 563955 358254
rect 563921 358220 563955 358234
rect 563921 358166 563955 358182
rect 563921 358148 563955 358166
rect 563921 358098 563955 358110
rect 563921 358076 563955 358098
rect 563921 358030 563955 358038
rect 563921 358004 563955 358030
rect 564179 358948 564213 358974
rect 564179 358940 564213 358948
rect 564179 358880 564213 358902
rect 564179 358868 564213 358880
rect 564179 358812 564213 358830
rect 564179 358796 564213 358812
rect 564179 358744 564213 358758
rect 564179 358724 564213 358744
rect 564179 358676 564213 358686
rect 564179 358652 564213 358676
rect 564179 358608 564213 358614
rect 564179 358580 564213 358608
rect 564179 358540 564213 358542
rect 564179 358508 564213 358540
rect 564179 358438 564213 358470
rect 564179 358436 564213 358438
rect 564179 358370 564213 358398
rect 564179 358364 564213 358370
rect 564179 358302 564213 358326
rect 564179 358292 564213 358302
rect 564179 358234 564213 358254
rect 564179 358220 564213 358234
rect 564179 358166 564213 358182
rect 564179 358148 564213 358166
rect 564179 358098 564213 358110
rect 564179 358076 564213 358098
rect 564179 358030 564213 358038
rect 564179 358004 564213 358030
rect 564437 358948 564471 358974
rect 564437 358940 564471 358948
rect 564437 358880 564471 358902
rect 564437 358868 564471 358880
rect 564437 358812 564471 358830
rect 564437 358796 564471 358812
rect 564437 358744 564471 358758
rect 564437 358724 564471 358744
rect 564437 358676 564471 358686
rect 564437 358652 564471 358676
rect 564437 358608 564471 358614
rect 564437 358580 564471 358608
rect 564437 358540 564471 358542
rect 564437 358508 564471 358540
rect 564437 358438 564471 358470
rect 564437 358436 564471 358438
rect 564437 358370 564471 358398
rect 564437 358364 564471 358370
rect 564437 358302 564471 358326
rect 564437 358292 564471 358302
rect 564437 358234 564471 358254
rect 564437 358220 564471 358234
rect 564437 358166 564471 358182
rect 564437 358148 564471 358166
rect 564437 358098 564471 358110
rect 564437 358076 564471 358098
rect 564437 358030 564471 358038
rect 564437 358004 564471 358030
rect 564695 358948 564729 358974
rect 564695 358940 564729 358948
rect 564695 358880 564729 358902
rect 564695 358868 564729 358880
rect 564695 358812 564729 358830
rect 564695 358796 564729 358812
rect 564695 358744 564729 358758
rect 564695 358724 564729 358744
rect 564695 358676 564729 358686
rect 564695 358652 564729 358676
rect 564695 358608 564729 358614
rect 564695 358580 564729 358608
rect 564695 358540 564729 358542
rect 564695 358508 564729 358540
rect 564695 358438 564729 358470
rect 564695 358436 564729 358438
rect 564695 358370 564729 358398
rect 564695 358364 564729 358370
rect 564695 358302 564729 358326
rect 564695 358292 564729 358302
rect 564695 358234 564729 358254
rect 564695 358220 564729 358234
rect 564695 358166 564729 358182
rect 564695 358148 564729 358166
rect 564695 358098 564729 358110
rect 564695 358076 564729 358098
rect 564695 358030 564729 358038
rect 564695 358004 564729 358030
rect 564953 358948 564987 358974
rect 564953 358940 564987 358948
rect 564953 358880 564987 358902
rect 564953 358868 564987 358880
rect 564953 358812 564987 358830
rect 564953 358796 564987 358812
rect 564953 358744 564987 358758
rect 564953 358724 564987 358744
rect 564953 358676 564987 358686
rect 564953 358652 564987 358676
rect 564953 358608 564987 358614
rect 564953 358580 564987 358608
rect 564953 358540 564987 358542
rect 564953 358508 564987 358540
rect 564953 358438 564987 358470
rect 564953 358436 564987 358438
rect 564953 358370 564987 358398
rect 564953 358364 564987 358370
rect 564953 358302 564987 358326
rect 564953 358292 564987 358302
rect 564953 358234 564987 358254
rect 564953 358220 564987 358234
rect 564953 358166 564987 358182
rect 564953 358148 564987 358166
rect 564953 358098 564987 358110
rect 564953 358076 564987 358098
rect 564953 358030 564987 358038
rect 564953 358004 564987 358030
rect 565211 358948 565245 358974
rect 565211 358940 565245 358948
rect 565211 358880 565245 358902
rect 565211 358868 565245 358880
rect 565211 358812 565245 358830
rect 565211 358796 565245 358812
rect 565211 358744 565245 358758
rect 565211 358724 565245 358744
rect 565211 358676 565245 358686
rect 565211 358652 565245 358676
rect 565211 358608 565245 358614
rect 565211 358580 565245 358608
rect 565211 358540 565245 358542
rect 565211 358508 565245 358540
rect 565211 358438 565245 358470
rect 565211 358436 565245 358438
rect 565211 358370 565245 358398
rect 565211 358364 565245 358370
rect 565211 358302 565245 358326
rect 565211 358292 565245 358302
rect 565211 358234 565245 358254
rect 565211 358220 565245 358234
rect 565211 358166 565245 358182
rect 565211 358148 565245 358166
rect 565211 358098 565245 358110
rect 565211 358076 565245 358098
rect 565211 358030 565245 358038
rect 565211 358004 565245 358030
rect 565469 358948 565503 358974
rect 565469 358940 565503 358948
rect 565469 358880 565503 358902
rect 565469 358868 565503 358880
rect 565469 358812 565503 358830
rect 565469 358796 565503 358812
rect 565469 358744 565503 358758
rect 565469 358724 565503 358744
rect 565469 358676 565503 358686
rect 565469 358652 565503 358676
rect 565469 358608 565503 358614
rect 565469 358580 565503 358608
rect 565469 358540 565503 358542
rect 565469 358508 565503 358540
rect 565469 358438 565503 358470
rect 565469 358436 565503 358438
rect 565469 358370 565503 358398
rect 565469 358364 565503 358370
rect 565469 358302 565503 358326
rect 565469 358292 565503 358302
rect 565469 358234 565503 358254
rect 565469 358220 565503 358234
rect 565469 358166 565503 358182
rect 565469 358148 565503 358166
rect 565469 358098 565503 358110
rect 565469 358076 565503 358098
rect 565469 358030 565503 358038
rect 565469 358004 565503 358030
rect 565727 358948 565761 358974
rect 565727 358940 565761 358948
rect 565727 358880 565761 358902
rect 565727 358868 565761 358880
rect 565727 358812 565761 358830
rect 565727 358796 565761 358812
rect 565727 358744 565761 358758
rect 565727 358724 565761 358744
rect 565727 358676 565761 358686
rect 565727 358652 565761 358676
rect 565727 358608 565761 358614
rect 565727 358580 565761 358608
rect 565727 358540 565761 358542
rect 565727 358508 565761 358540
rect 565727 358438 565761 358470
rect 565727 358436 565761 358438
rect 565727 358370 565761 358398
rect 565727 358364 565761 358370
rect 565727 358302 565761 358326
rect 565727 358292 565761 358302
rect 565727 358234 565761 358254
rect 565727 358220 565761 358234
rect 565727 358166 565761 358182
rect 565727 358148 565761 358166
rect 565727 358098 565761 358110
rect 565727 358076 565761 358098
rect 565727 358030 565761 358038
rect 565727 358004 565761 358030
rect 566007 357870 566113 357976
rect 574705 358878 574739 358904
rect 574705 358870 574739 358878
rect 574705 358810 574739 358832
rect 574705 358798 574739 358810
rect 574705 358742 574739 358760
rect 574705 358726 574739 358742
rect 574705 358674 574739 358688
rect 574705 358654 574739 358674
rect 574705 358606 574739 358616
rect 574705 358582 574739 358606
rect 574705 358538 574739 358544
rect 574705 358510 574739 358538
rect 574705 358470 574739 358472
rect 574705 358438 574739 358470
rect 574705 358368 574739 358400
rect 574705 358366 574739 358368
rect 574705 358300 574739 358328
rect 574705 358294 574739 358300
rect 574705 358232 574739 358256
rect 574705 358222 574739 358232
rect 574705 358164 574739 358184
rect 574705 358150 574739 358164
rect 574705 358096 574739 358112
rect 574705 358078 574739 358096
rect 574705 358028 574739 358040
rect 574705 358006 574739 358028
rect 574705 357960 574739 357968
rect 574705 357934 574739 357960
rect 574963 358878 574997 358904
rect 574963 358870 574997 358878
rect 574963 358810 574997 358832
rect 574963 358798 574997 358810
rect 574963 358742 574997 358760
rect 574963 358726 574997 358742
rect 574963 358674 574997 358688
rect 574963 358654 574997 358674
rect 574963 358606 574997 358616
rect 574963 358582 574997 358606
rect 574963 358538 574997 358544
rect 574963 358510 574997 358538
rect 574963 358470 574997 358472
rect 574963 358438 574997 358470
rect 574963 358368 574997 358400
rect 574963 358366 574997 358368
rect 574963 358300 574997 358328
rect 574963 358294 574997 358300
rect 574963 358232 574997 358256
rect 574963 358222 574997 358232
rect 574963 358164 574997 358184
rect 574963 358150 574997 358164
rect 574963 358096 574997 358112
rect 574963 358078 574997 358096
rect 574963 358028 574997 358040
rect 574963 358006 574997 358028
rect 574963 357960 574997 357968
rect 574963 357934 574997 357960
rect 575221 358878 575255 358904
rect 575221 358870 575255 358878
rect 575221 358810 575255 358832
rect 575221 358798 575255 358810
rect 575221 358742 575255 358760
rect 575221 358726 575255 358742
rect 575221 358674 575255 358688
rect 575221 358654 575255 358674
rect 575221 358606 575255 358616
rect 575221 358582 575255 358606
rect 575221 358538 575255 358544
rect 575221 358510 575255 358538
rect 575221 358470 575255 358472
rect 575221 358438 575255 358470
rect 575221 358368 575255 358400
rect 575221 358366 575255 358368
rect 575221 358300 575255 358328
rect 575221 358294 575255 358300
rect 575221 358232 575255 358256
rect 575221 358222 575255 358232
rect 575221 358164 575255 358184
rect 575221 358150 575255 358164
rect 575221 358096 575255 358112
rect 575221 358078 575255 358096
rect 575221 358028 575255 358040
rect 575221 358006 575255 358028
rect 575221 357960 575255 357968
rect 575221 357934 575255 357960
rect 575479 358878 575513 358904
rect 575479 358870 575513 358878
rect 575479 358810 575513 358832
rect 575479 358798 575513 358810
rect 575479 358742 575513 358760
rect 575479 358726 575513 358742
rect 575479 358674 575513 358688
rect 575479 358654 575513 358674
rect 575479 358606 575513 358616
rect 575479 358582 575513 358606
rect 575479 358538 575513 358544
rect 575479 358510 575513 358538
rect 575479 358470 575513 358472
rect 575479 358438 575513 358470
rect 575479 358368 575513 358400
rect 575479 358366 575513 358368
rect 575479 358300 575513 358328
rect 575479 358294 575513 358300
rect 575479 358232 575513 358256
rect 575479 358222 575513 358232
rect 575479 358164 575513 358184
rect 575479 358150 575513 358164
rect 575479 358096 575513 358112
rect 575479 358078 575513 358096
rect 575479 358028 575513 358040
rect 575479 358006 575513 358028
rect 575479 357960 575513 357968
rect 575479 357934 575513 357960
rect 575737 358878 575771 358904
rect 575737 358870 575771 358878
rect 575737 358810 575771 358832
rect 575737 358798 575771 358810
rect 575737 358742 575771 358760
rect 575737 358726 575771 358742
rect 575737 358674 575771 358688
rect 575737 358654 575771 358674
rect 575737 358606 575771 358616
rect 575737 358582 575771 358606
rect 575737 358538 575771 358544
rect 575737 358510 575771 358538
rect 575737 358470 575771 358472
rect 575737 358438 575771 358470
rect 575737 358368 575771 358400
rect 575737 358366 575771 358368
rect 575737 358300 575771 358328
rect 575737 358294 575771 358300
rect 575737 358232 575771 358256
rect 575737 358222 575771 358232
rect 575737 358164 575771 358184
rect 575737 358150 575771 358164
rect 575737 358096 575771 358112
rect 575737 358078 575771 358096
rect 575737 358028 575771 358040
rect 575737 358006 575771 358028
rect 575737 357960 575771 357968
rect 575737 357934 575771 357960
rect 575995 358878 576029 358904
rect 575995 358870 576029 358878
rect 575995 358810 576029 358832
rect 575995 358798 576029 358810
rect 575995 358742 576029 358760
rect 575995 358726 576029 358742
rect 575995 358674 576029 358688
rect 575995 358654 576029 358674
rect 575995 358606 576029 358616
rect 575995 358582 576029 358606
rect 575995 358538 576029 358544
rect 575995 358510 576029 358538
rect 575995 358470 576029 358472
rect 575995 358438 576029 358470
rect 575995 358368 576029 358400
rect 575995 358366 576029 358368
rect 575995 358300 576029 358328
rect 575995 358294 576029 358300
rect 575995 358232 576029 358256
rect 575995 358222 576029 358232
rect 575995 358164 576029 358184
rect 575995 358150 576029 358164
rect 575995 358096 576029 358112
rect 575995 358078 576029 358096
rect 575995 358028 576029 358040
rect 575995 358006 576029 358028
rect 575995 357960 576029 357968
rect 575995 357934 576029 357960
rect 576253 358878 576287 358904
rect 576253 358870 576287 358878
rect 576253 358810 576287 358832
rect 576253 358798 576287 358810
rect 576253 358742 576287 358760
rect 576253 358726 576287 358742
rect 576253 358674 576287 358688
rect 576253 358654 576287 358674
rect 576253 358606 576287 358616
rect 576253 358582 576287 358606
rect 576253 358538 576287 358544
rect 576253 358510 576287 358538
rect 576253 358470 576287 358472
rect 576253 358438 576287 358470
rect 576253 358368 576287 358400
rect 576253 358366 576287 358368
rect 576253 358300 576287 358328
rect 576253 358294 576287 358300
rect 576253 358232 576287 358256
rect 576253 358222 576287 358232
rect 576253 358164 576287 358184
rect 576253 358150 576287 358164
rect 576253 358096 576287 358112
rect 576253 358078 576287 358096
rect 576253 358028 576287 358040
rect 576253 358006 576287 358028
rect 576253 357960 576287 357968
rect 576253 357934 576287 357960
rect 576511 358878 576545 358904
rect 576511 358870 576545 358878
rect 576511 358810 576545 358832
rect 576511 358798 576545 358810
rect 576511 358742 576545 358760
rect 576511 358726 576545 358742
rect 576511 358674 576545 358688
rect 576511 358654 576545 358674
rect 576511 358606 576545 358616
rect 576511 358582 576545 358606
rect 576511 358538 576545 358544
rect 576511 358510 576545 358538
rect 576511 358470 576545 358472
rect 576511 358438 576545 358470
rect 576511 358368 576545 358400
rect 576511 358366 576545 358368
rect 576511 358300 576545 358328
rect 576511 358294 576545 358300
rect 576511 358232 576545 358256
rect 576511 358222 576545 358232
rect 576511 358164 576545 358184
rect 576511 358150 576545 358164
rect 576511 358096 576545 358112
rect 576511 358078 576545 358096
rect 576511 358028 576545 358040
rect 576511 358006 576545 358028
rect 576511 357960 576545 357968
rect 576511 357934 576545 357960
rect 576769 358878 576803 358904
rect 576769 358870 576803 358878
rect 576769 358810 576803 358832
rect 576769 358798 576803 358810
rect 576769 358742 576803 358760
rect 576769 358726 576803 358742
rect 576769 358674 576803 358688
rect 576769 358654 576803 358674
rect 576769 358606 576803 358616
rect 576769 358582 576803 358606
rect 576769 358538 576803 358544
rect 576769 358510 576803 358538
rect 576769 358470 576803 358472
rect 576769 358438 576803 358470
rect 576769 358368 576803 358400
rect 576769 358366 576803 358368
rect 576769 358300 576803 358328
rect 576769 358294 576803 358300
rect 576769 358232 576803 358256
rect 576769 358222 576803 358232
rect 576769 358164 576803 358184
rect 576769 358150 576803 358164
rect 576769 358096 576803 358112
rect 576769 358078 576803 358096
rect 576769 358028 576803 358040
rect 576769 358006 576803 358028
rect 576769 357960 576803 357968
rect 576769 357934 576803 357960
rect 577027 358878 577061 358904
rect 577027 358870 577061 358878
rect 577027 358810 577061 358832
rect 577027 358798 577061 358810
rect 577027 358742 577061 358760
rect 577027 358726 577061 358742
rect 577027 358674 577061 358688
rect 577027 358654 577061 358674
rect 577027 358606 577061 358616
rect 577027 358582 577061 358606
rect 577027 358538 577061 358544
rect 577027 358510 577061 358538
rect 577027 358470 577061 358472
rect 577027 358438 577061 358470
rect 577027 358368 577061 358400
rect 577027 358366 577061 358368
rect 577027 358300 577061 358328
rect 577027 358294 577061 358300
rect 577027 358232 577061 358256
rect 577027 358222 577061 358232
rect 577027 358164 577061 358184
rect 577027 358150 577061 358164
rect 577027 358096 577061 358112
rect 577027 358078 577061 358096
rect 577027 358028 577061 358040
rect 577027 358006 577061 358028
rect 577027 357960 577061 357968
rect 577027 357934 577061 357960
rect 577285 358878 577319 358904
rect 577285 358870 577319 358878
rect 577285 358810 577319 358832
rect 577285 358798 577319 358810
rect 577285 358742 577319 358760
rect 577285 358726 577319 358742
rect 577285 358674 577319 358688
rect 577285 358654 577319 358674
rect 577285 358606 577319 358616
rect 577285 358582 577319 358606
rect 577285 358538 577319 358544
rect 577285 358510 577319 358538
rect 577285 358470 577319 358472
rect 577285 358438 577319 358470
rect 577285 358368 577319 358400
rect 577285 358366 577319 358368
rect 577285 358300 577319 358328
rect 577285 358294 577319 358300
rect 577285 358232 577319 358256
rect 577285 358222 577319 358232
rect 577285 358164 577319 358184
rect 577285 358150 577319 358164
rect 577285 358096 577319 358112
rect 577285 358078 577319 358096
rect 577285 358028 577319 358040
rect 577285 358006 577319 358028
rect 577285 357960 577319 357968
rect 577285 357934 577319 357960
rect 577543 358878 577577 358904
rect 577543 358870 577577 358878
rect 577543 358810 577577 358832
rect 577543 358798 577577 358810
rect 577543 358742 577577 358760
rect 577543 358726 577577 358742
rect 577543 358674 577577 358688
rect 577543 358654 577577 358674
rect 577543 358606 577577 358616
rect 577543 358582 577577 358606
rect 577543 358538 577577 358544
rect 577543 358510 577577 358538
rect 577543 358470 577577 358472
rect 577543 358438 577577 358470
rect 577543 358368 577577 358400
rect 577543 358366 577577 358368
rect 577543 358300 577577 358328
rect 577543 358294 577577 358300
rect 577543 358232 577577 358256
rect 577543 358222 577577 358232
rect 577543 358164 577577 358184
rect 577543 358150 577577 358164
rect 577543 358096 577577 358112
rect 577543 358078 577577 358096
rect 577543 358028 577577 358040
rect 577543 358006 577577 358028
rect 577543 357960 577577 357968
rect 577543 357934 577577 357960
rect 577801 358878 577835 358904
rect 577801 358870 577835 358878
rect 577801 358810 577835 358832
rect 577801 358798 577835 358810
rect 577801 358742 577835 358760
rect 577801 358726 577835 358742
rect 577801 358674 577835 358688
rect 577801 358654 577835 358674
rect 577801 358606 577835 358616
rect 577801 358582 577835 358606
rect 577801 358538 577835 358544
rect 577801 358510 577835 358538
rect 577801 358470 577835 358472
rect 577801 358438 577835 358470
rect 577801 358368 577835 358400
rect 577801 358366 577835 358368
rect 577801 358300 577835 358328
rect 577801 358294 577835 358300
rect 577801 358232 577835 358256
rect 577801 358222 577835 358232
rect 577801 358164 577835 358184
rect 577801 358150 577835 358164
rect 577801 358096 577835 358112
rect 577801 358078 577835 358096
rect 577801 358028 577835 358040
rect 577801 358006 577835 358028
rect 577801 357960 577835 357968
rect 577801 357934 577835 357960
rect 578059 358878 578093 358904
rect 578059 358870 578093 358878
rect 578059 358810 578093 358832
rect 578059 358798 578093 358810
rect 578059 358742 578093 358760
rect 578059 358726 578093 358742
rect 578059 358674 578093 358688
rect 578059 358654 578093 358674
rect 578059 358606 578093 358616
rect 578059 358582 578093 358606
rect 578059 358538 578093 358544
rect 578059 358510 578093 358538
rect 578059 358470 578093 358472
rect 578059 358438 578093 358470
rect 578059 358368 578093 358400
rect 578059 358366 578093 358368
rect 578059 358300 578093 358328
rect 578059 358294 578093 358300
rect 578059 358232 578093 358256
rect 578059 358222 578093 358232
rect 578059 358164 578093 358184
rect 578059 358150 578093 358164
rect 578059 358096 578093 358112
rect 578059 358078 578093 358096
rect 578059 358028 578093 358040
rect 578059 358006 578093 358028
rect 578059 357960 578093 357968
rect 578059 357934 578093 357960
rect 578317 358878 578351 358904
rect 578317 358870 578351 358878
rect 578317 358810 578351 358832
rect 578317 358798 578351 358810
rect 578317 358742 578351 358760
rect 578317 358726 578351 358742
rect 578317 358674 578351 358688
rect 578317 358654 578351 358674
rect 578317 358606 578351 358616
rect 578317 358582 578351 358606
rect 578317 358538 578351 358544
rect 578317 358510 578351 358538
rect 578317 358470 578351 358472
rect 578317 358438 578351 358470
rect 578317 358368 578351 358400
rect 578317 358366 578351 358368
rect 578317 358300 578351 358328
rect 578317 358294 578351 358300
rect 578317 358232 578351 358256
rect 578317 358222 578351 358232
rect 578317 358164 578351 358184
rect 578317 358150 578351 358164
rect 578317 358096 578351 358112
rect 578317 358078 578351 358096
rect 578317 358028 578351 358040
rect 578317 358006 578351 358028
rect 578317 357960 578351 357968
rect 578317 357934 578351 357960
rect 578575 358878 578609 358904
rect 578575 358870 578609 358878
rect 578575 358810 578609 358832
rect 578575 358798 578609 358810
rect 578575 358742 578609 358760
rect 578575 358726 578609 358742
rect 578575 358674 578609 358688
rect 578575 358654 578609 358674
rect 578575 358606 578609 358616
rect 578575 358582 578609 358606
rect 578575 358538 578609 358544
rect 578575 358510 578609 358538
rect 578575 358470 578609 358472
rect 578575 358438 578609 358470
rect 578575 358368 578609 358400
rect 578575 358366 578609 358368
rect 578575 358300 578609 358328
rect 578575 358294 578609 358300
rect 578575 358232 578609 358256
rect 578575 358222 578609 358232
rect 578575 358164 578609 358184
rect 578575 358150 578609 358164
rect 578575 358096 578609 358112
rect 578575 358078 578609 358096
rect 578575 358028 578609 358040
rect 578575 358006 578609 358028
rect 578575 357960 578609 357968
rect 578575 357934 578609 357960
rect 578833 358878 578867 358904
rect 578833 358870 578867 358878
rect 578833 358810 578867 358832
rect 578833 358798 578867 358810
rect 578833 358742 578867 358760
rect 578833 358726 578867 358742
rect 578833 358674 578867 358688
rect 578833 358654 578867 358674
rect 578833 358606 578867 358616
rect 578833 358582 578867 358606
rect 578833 358538 578867 358544
rect 578833 358510 578867 358538
rect 578833 358470 578867 358472
rect 578833 358438 578867 358470
rect 578833 358368 578867 358400
rect 578833 358366 578867 358368
rect 578833 358300 578867 358328
rect 578833 358294 578867 358300
rect 578833 358232 578867 358256
rect 578833 358222 578867 358232
rect 578833 358164 578867 358184
rect 578833 358150 578867 358164
rect 578833 358096 578867 358112
rect 578833 358078 578867 358096
rect 578833 358028 578867 358040
rect 578833 358006 578867 358028
rect 578833 357960 578867 357968
rect 578833 357934 578867 357960
rect 579091 358878 579125 358904
rect 579091 358870 579125 358878
rect 579091 358810 579125 358832
rect 579091 358798 579125 358810
rect 579091 358742 579125 358760
rect 579091 358726 579125 358742
rect 579091 358674 579125 358688
rect 579091 358654 579125 358674
rect 579091 358606 579125 358616
rect 579091 358582 579125 358606
rect 579091 358538 579125 358544
rect 579091 358510 579125 358538
rect 579091 358470 579125 358472
rect 579091 358438 579125 358470
rect 579091 358368 579125 358400
rect 579091 358366 579125 358368
rect 579091 358300 579125 358328
rect 579091 358294 579125 358300
rect 579091 358232 579125 358256
rect 579091 358222 579125 358232
rect 579091 358164 579125 358184
rect 579091 358150 579125 358164
rect 579091 358096 579125 358112
rect 579091 358078 579125 358096
rect 579091 358028 579125 358040
rect 579091 358006 579125 358028
rect 579091 357960 579125 357968
rect 579091 357934 579125 357960
rect 579349 358878 579383 358904
rect 579349 358870 579383 358878
rect 579349 358810 579383 358832
rect 579349 358798 579383 358810
rect 579349 358742 579383 358760
rect 579349 358726 579383 358742
rect 579349 358674 579383 358688
rect 579349 358654 579383 358674
rect 579349 358606 579383 358616
rect 579349 358582 579383 358606
rect 579349 358538 579383 358544
rect 579349 358510 579383 358538
rect 579349 358470 579383 358472
rect 579349 358438 579383 358470
rect 579349 358368 579383 358400
rect 579349 358366 579383 358368
rect 579349 358300 579383 358328
rect 579349 358294 579383 358300
rect 579349 358232 579383 358256
rect 579349 358222 579383 358232
rect 579349 358164 579383 358184
rect 579349 358150 579383 358164
rect 579349 358096 579383 358112
rect 579349 358078 579383 358096
rect 579349 358028 579383 358040
rect 579349 358006 579383 358028
rect 579349 357960 579383 357968
rect 579349 357934 579383 357960
rect 579607 358878 579641 358904
rect 579607 358870 579641 358878
rect 579607 358810 579641 358832
rect 579607 358798 579641 358810
rect 579607 358742 579641 358760
rect 579607 358726 579641 358742
rect 579607 358674 579641 358688
rect 579607 358654 579641 358674
rect 579607 358606 579641 358616
rect 579607 358582 579641 358606
rect 579607 358538 579641 358544
rect 579607 358510 579641 358538
rect 579607 358470 579641 358472
rect 579607 358438 579641 358470
rect 579607 358368 579641 358400
rect 579607 358366 579641 358368
rect 579607 358300 579641 358328
rect 579607 358294 579641 358300
rect 579607 358232 579641 358256
rect 579607 358222 579641 358232
rect 579607 358164 579641 358184
rect 579607 358150 579641 358164
rect 579607 358096 579641 358112
rect 579607 358078 579641 358096
rect 579607 358028 579641 358040
rect 579607 358006 579641 358028
rect 579607 357960 579641 357968
rect 579607 357934 579641 357960
rect 579865 358878 579899 358904
rect 579865 358870 579899 358878
rect 579865 358810 579899 358832
rect 579865 358798 579899 358810
rect 579865 358742 579899 358760
rect 579865 358726 579899 358742
rect 579865 358674 579899 358688
rect 579865 358654 579899 358674
rect 579865 358606 579899 358616
rect 579865 358582 579899 358606
rect 579865 358538 579899 358544
rect 579865 358510 579899 358538
rect 579865 358470 579899 358472
rect 579865 358438 579899 358470
rect 579865 358368 579899 358400
rect 579865 358366 579899 358368
rect 579865 358300 579899 358328
rect 579865 358294 579899 358300
rect 579865 358232 579899 358256
rect 579865 358222 579899 358232
rect 579865 358164 579899 358184
rect 579865 358150 579899 358164
rect 579865 358096 579899 358112
rect 579865 358078 579899 358096
rect 579865 358028 579899 358040
rect 579865 358006 579899 358028
rect 579865 357960 579899 357968
rect 579865 357934 579899 357960
rect 580058 357762 580092 357796
rect 574451 357620 574485 357654
rect 560755 357472 560789 357506
rect 560955 357472 560989 357506
rect 561155 357472 561189 357506
rect 561355 357472 561389 357506
rect 561555 357472 561589 357506
rect 561755 357472 561789 357506
rect 561955 357472 561989 357506
rect 562155 357472 562189 357506
rect 562355 357472 562389 357506
rect 562555 357472 562589 357506
rect 562755 357472 562789 357506
rect 562955 357472 562989 357506
rect 563155 357472 563189 357506
rect 563355 357472 563389 357506
rect 563555 357472 563589 357506
rect 563755 357472 563789 357506
rect 563955 357472 563989 357506
rect 564155 357472 564189 357506
rect 564355 357472 564389 357506
rect 564555 357472 564589 357506
rect 564755 357472 564789 357506
rect 564955 357472 564989 357506
rect 565155 357472 565189 357506
rect 565355 357472 565389 357506
rect 565555 357472 565589 357506
rect 574729 357402 574763 357436
rect 574929 357402 574963 357436
rect 575129 357402 575163 357436
rect 575329 357402 575363 357436
rect 575529 357402 575563 357436
rect 575729 357402 575763 357436
rect 575929 357402 575963 357436
rect 576129 357402 576163 357436
rect 576329 357402 576363 357436
rect 576529 357402 576563 357436
rect 576729 357402 576763 357436
rect 576929 357402 576963 357436
rect 577129 357402 577163 357436
rect 577329 357402 577363 357436
rect 577529 357402 577563 357436
rect 577729 357402 577763 357436
rect 577929 357402 577963 357436
rect 578129 357402 578163 357436
rect 578329 357402 578363 357436
rect 578529 357402 578563 357436
rect 578729 357402 578763 357436
rect 578929 357402 578963 357436
rect 579129 357402 579163 357436
rect 579329 357402 579363 357436
rect 579529 357402 579563 357436
rect 579729 357402 579763 357436
rect 575177 313114 575211 313148
rect 575377 313114 575411 313148
rect 575577 313114 575611 313148
rect 575777 313114 575811 313148
rect 575977 313114 576011 313148
rect 576177 313114 576211 313148
rect 576377 313114 576411 313148
rect 576577 313114 576611 313148
rect 576777 313114 576811 313148
rect 576977 313114 577011 313148
rect 577177 313114 577211 313148
rect 577377 313114 577411 313148
rect 577577 313114 577611 313148
rect 577777 313114 577811 313148
rect 577977 313114 578011 313148
rect 578177 313114 578211 313148
rect 578377 313114 578411 313148
rect 578577 313114 578611 313148
rect 578777 313114 578811 313148
rect 578977 313114 579011 313148
rect 579177 313114 579211 313148
rect 579377 313114 579411 313148
rect 579577 313114 579611 313148
rect 579777 313114 579811 313148
rect 579977 313114 580011 313148
rect 580177 313114 580211 313148
rect 560617 313044 560651 313078
rect 560817 313044 560851 313078
rect 561017 313044 561051 313078
rect 561217 313044 561251 313078
rect 561417 313044 561451 313078
rect 561617 313044 561651 313078
rect 561817 313044 561851 313078
rect 562017 313044 562051 313078
rect 562217 313044 562251 313078
rect 562417 313044 562451 313078
rect 562617 313044 562651 313078
rect 562817 313044 562851 313078
rect 563017 313044 563051 313078
rect 563217 313044 563251 313078
rect 563417 313044 563451 313078
rect 563617 313044 563651 313078
rect 563817 313044 563851 313078
rect 564017 313044 564051 313078
rect 564217 313044 564251 313078
rect 564417 313044 564451 313078
rect 564617 313044 564651 313078
rect 564817 313044 564851 313078
rect 565017 313044 565051 313078
rect 565217 313044 565251 313078
rect 565417 313044 565451 313078
rect 560121 311595 560227 311701
rect 560429 312640 560463 312666
rect 560429 312632 560463 312640
rect 560429 312572 560463 312594
rect 560429 312560 560463 312572
rect 560429 312504 560463 312522
rect 560429 312488 560463 312504
rect 560429 312436 560463 312450
rect 560429 312416 560463 312436
rect 560429 312368 560463 312378
rect 560429 312344 560463 312368
rect 560429 312300 560463 312306
rect 560429 312272 560463 312300
rect 560429 312232 560463 312234
rect 560429 312200 560463 312232
rect 560429 312130 560463 312162
rect 560429 312128 560463 312130
rect 560429 312062 560463 312090
rect 560429 312056 560463 312062
rect 560429 311994 560463 312018
rect 560429 311984 560463 311994
rect 560429 311926 560463 311946
rect 560429 311912 560463 311926
rect 560429 311858 560463 311874
rect 560429 311840 560463 311858
rect 560429 311790 560463 311802
rect 560429 311768 560463 311790
rect 560429 311722 560463 311730
rect 560429 311696 560463 311722
rect 560687 312640 560721 312666
rect 560687 312632 560721 312640
rect 560687 312572 560721 312594
rect 560687 312560 560721 312572
rect 560687 312504 560721 312522
rect 560687 312488 560721 312504
rect 560687 312436 560721 312450
rect 560687 312416 560721 312436
rect 560687 312368 560721 312378
rect 560687 312344 560721 312368
rect 560687 312300 560721 312306
rect 560687 312272 560721 312300
rect 560687 312232 560721 312234
rect 560687 312200 560721 312232
rect 560687 312130 560721 312162
rect 560687 312128 560721 312130
rect 560687 312062 560721 312090
rect 560687 312056 560721 312062
rect 560687 311994 560721 312018
rect 560687 311984 560721 311994
rect 560687 311926 560721 311946
rect 560687 311912 560721 311926
rect 560687 311858 560721 311874
rect 560687 311840 560721 311858
rect 560687 311790 560721 311802
rect 560687 311768 560721 311790
rect 560687 311722 560721 311730
rect 560687 311696 560721 311722
rect 560945 312640 560979 312666
rect 560945 312632 560979 312640
rect 560945 312572 560979 312594
rect 560945 312560 560979 312572
rect 560945 312504 560979 312522
rect 560945 312488 560979 312504
rect 560945 312436 560979 312450
rect 560945 312416 560979 312436
rect 560945 312368 560979 312378
rect 560945 312344 560979 312368
rect 560945 312300 560979 312306
rect 560945 312272 560979 312300
rect 560945 312232 560979 312234
rect 560945 312200 560979 312232
rect 560945 312130 560979 312162
rect 560945 312128 560979 312130
rect 560945 312062 560979 312090
rect 560945 312056 560979 312062
rect 560945 311994 560979 312018
rect 560945 311984 560979 311994
rect 560945 311926 560979 311946
rect 560945 311912 560979 311926
rect 560945 311858 560979 311874
rect 560945 311840 560979 311858
rect 560945 311790 560979 311802
rect 560945 311768 560979 311790
rect 560945 311722 560979 311730
rect 560945 311696 560979 311722
rect 561203 312640 561237 312666
rect 561203 312632 561237 312640
rect 561203 312572 561237 312594
rect 561203 312560 561237 312572
rect 561203 312504 561237 312522
rect 561203 312488 561237 312504
rect 561203 312436 561237 312450
rect 561203 312416 561237 312436
rect 561203 312368 561237 312378
rect 561203 312344 561237 312368
rect 561203 312300 561237 312306
rect 561203 312272 561237 312300
rect 561203 312232 561237 312234
rect 561203 312200 561237 312232
rect 561203 312130 561237 312162
rect 561203 312128 561237 312130
rect 561203 312062 561237 312090
rect 561203 312056 561237 312062
rect 561203 311994 561237 312018
rect 561203 311984 561237 311994
rect 561203 311926 561237 311946
rect 561203 311912 561237 311926
rect 561203 311858 561237 311874
rect 561203 311840 561237 311858
rect 561203 311790 561237 311802
rect 561203 311768 561237 311790
rect 561203 311722 561237 311730
rect 561203 311696 561237 311722
rect 561461 312640 561495 312666
rect 561461 312632 561495 312640
rect 561461 312572 561495 312594
rect 561461 312560 561495 312572
rect 561461 312504 561495 312522
rect 561461 312488 561495 312504
rect 561461 312436 561495 312450
rect 561461 312416 561495 312436
rect 561461 312368 561495 312378
rect 561461 312344 561495 312368
rect 561461 312300 561495 312306
rect 561461 312272 561495 312300
rect 561461 312232 561495 312234
rect 561461 312200 561495 312232
rect 561461 312130 561495 312162
rect 561461 312128 561495 312130
rect 561461 312062 561495 312090
rect 561461 312056 561495 312062
rect 561461 311994 561495 312018
rect 561461 311984 561495 311994
rect 561461 311926 561495 311946
rect 561461 311912 561495 311926
rect 561461 311858 561495 311874
rect 561461 311840 561495 311858
rect 561461 311790 561495 311802
rect 561461 311768 561495 311790
rect 561461 311722 561495 311730
rect 561461 311696 561495 311722
rect 561719 312640 561753 312666
rect 561719 312632 561753 312640
rect 561719 312572 561753 312594
rect 561719 312560 561753 312572
rect 561719 312504 561753 312522
rect 561719 312488 561753 312504
rect 561719 312436 561753 312450
rect 561719 312416 561753 312436
rect 561719 312368 561753 312378
rect 561719 312344 561753 312368
rect 561719 312300 561753 312306
rect 561719 312272 561753 312300
rect 561719 312232 561753 312234
rect 561719 312200 561753 312232
rect 561719 312130 561753 312162
rect 561719 312128 561753 312130
rect 561719 312062 561753 312090
rect 561719 312056 561753 312062
rect 561719 311994 561753 312018
rect 561719 311984 561753 311994
rect 561719 311926 561753 311946
rect 561719 311912 561753 311926
rect 561719 311858 561753 311874
rect 561719 311840 561753 311858
rect 561719 311790 561753 311802
rect 561719 311768 561753 311790
rect 561719 311722 561753 311730
rect 561719 311696 561753 311722
rect 561977 312640 562011 312666
rect 561977 312632 562011 312640
rect 561977 312572 562011 312594
rect 561977 312560 562011 312572
rect 561977 312504 562011 312522
rect 561977 312488 562011 312504
rect 561977 312436 562011 312450
rect 561977 312416 562011 312436
rect 561977 312368 562011 312378
rect 561977 312344 562011 312368
rect 561977 312300 562011 312306
rect 561977 312272 562011 312300
rect 561977 312232 562011 312234
rect 561977 312200 562011 312232
rect 561977 312130 562011 312162
rect 561977 312128 562011 312130
rect 561977 312062 562011 312090
rect 561977 312056 562011 312062
rect 561977 311994 562011 312018
rect 561977 311984 562011 311994
rect 561977 311926 562011 311946
rect 561977 311912 562011 311926
rect 561977 311858 562011 311874
rect 561977 311840 562011 311858
rect 561977 311790 562011 311802
rect 561977 311768 562011 311790
rect 561977 311722 562011 311730
rect 561977 311696 562011 311722
rect 562235 312640 562269 312666
rect 562235 312632 562269 312640
rect 562235 312572 562269 312594
rect 562235 312560 562269 312572
rect 562235 312504 562269 312522
rect 562235 312488 562269 312504
rect 562235 312436 562269 312450
rect 562235 312416 562269 312436
rect 562235 312368 562269 312378
rect 562235 312344 562269 312368
rect 562235 312300 562269 312306
rect 562235 312272 562269 312300
rect 562235 312232 562269 312234
rect 562235 312200 562269 312232
rect 562235 312130 562269 312162
rect 562235 312128 562269 312130
rect 562235 312062 562269 312090
rect 562235 312056 562269 312062
rect 562235 311994 562269 312018
rect 562235 311984 562269 311994
rect 562235 311926 562269 311946
rect 562235 311912 562269 311926
rect 562235 311858 562269 311874
rect 562235 311840 562269 311858
rect 562235 311790 562269 311802
rect 562235 311768 562269 311790
rect 562235 311722 562269 311730
rect 562235 311696 562269 311722
rect 562493 312640 562527 312666
rect 562493 312632 562527 312640
rect 562493 312572 562527 312594
rect 562493 312560 562527 312572
rect 562493 312504 562527 312522
rect 562493 312488 562527 312504
rect 562493 312436 562527 312450
rect 562493 312416 562527 312436
rect 562493 312368 562527 312378
rect 562493 312344 562527 312368
rect 562493 312300 562527 312306
rect 562493 312272 562527 312300
rect 562493 312232 562527 312234
rect 562493 312200 562527 312232
rect 562493 312130 562527 312162
rect 562493 312128 562527 312130
rect 562493 312062 562527 312090
rect 562493 312056 562527 312062
rect 562493 311994 562527 312018
rect 562493 311984 562527 311994
rect 562493 311926 562527 311946
rect 562493 311912 562527 311926
rect 562493 311858 562527 311874
rect 562493 311840 562527 311858
rect 562493 311790 562527 311802
rect 562493 311768 562527 311790
rect 562493 311722 562527 311730
rect 562493 311696 562527 311722
rect 562751 312640 562785 312666
rect 562751 312632 562785 312640
rect 562751 312572 562785 312594
rect 562751 312560 562785 312572
rect 562751 312504 562785 312522
rect 562751 312488 562785 312504
rect 562751 312436 562785 312450
rect 562751 312416 562785 312436
rect 562751 312368 562785 312378
rect 562751 312344 562785 312368
rect 562751 312300 562785 312306
rect 562751 312272 562785 312300
rect 562751 312232 562785 312234
rect 562751 312200 562785 312232
rect 562751 312130 562785 312162
rect 562751 312128 562785 312130
rect 562751 312062 562785 312090
rect 562751 312056 562785 312062
rect 562751 311994 562785 312018
rect 562751 311984 562785 311994
rect 562751 311926 562785 311946
rect 562751 311912 562785 311926
rect 562751 311858 562785 311874
rect 562751 311840 562785 311858
rect 562751 311790 562785 311802
rect 562751 311768 562785 311790
rect 562751 311722 562785 311730
rect 562751 311696 562785 311722
rect 563009 312640 563043 312666
rect 563009 312632 563043 312640
rect 563009 312572 563043 312594
rect 563009 312560 563043 312572
rect 563009 312504 563043 312522
rect 563009 312488 563043 312504
rect 563009 312436 563043 312450
rect 563009 312416 563043 312436
rect 563009 312368 563043 312378
rect 563009 312344 563043 312368
rect 563009 312300 563043 312306
rect 563009 312272 563043 312300
rect 563009 312232 563043 312234
rect 563009 312200 563043 312232
rect 563009 312130 563043 312162
rect 563009 312128 563043 312130
rect 563009 312062 563043 312090
rect 563009 312056 563043 312062
rect 563009 311994 563043 312018
rect 563009 311984 563043 311994
rect 563009 311926 563043 311946
rect 563009 311912 563043 311926
rect 563009 311858 563043 311874
rect 563009 311840 563043 311858
rect 563009 311790 563043 311802
rect 563009 311768 563043 311790
rect 563009 311722 563043 311730
rect 563009 311696 563043 311722
rect 563267 312640 563301 312666
rect 563267 312632 563301 312640
rect 563267 312572 563301 312594
rect 563267 312560 563301 312572
rect 563267 312504 563301 312522
rect 563267 312488 563301 312504
rect 563267 312436 563301 312450
rect 563267 312416 563301 312436
rect 563267 312368 563301 312378
rect 563267 312344 563301 312368
rect 563267 312300 563301 312306
rect 563267 312272 563301 312300
rect 563267 312232 563301 312234
rect 563267 312200 563301 312232
rect 563267 312130 563301 312162
rect 563267 312128 563301 312130
rect 563267 312062 563301 312090
rect 563267 312056 563301 312062
rect 563267 311994 563301 312018
rect 563267 311984 563301 311994
rect 563267 311926 563301 311946
rect 563267 311912 563301 311926
rect 563267 311858 563301 311874
rect 563267 311840 563301 311858
rect 563267 311790 563301 311802
rect 563267 311768 563301 311790
rect 563267 311722 563301 311730
rect 563267 311696 563301 311722
rect 563525 312640 563559 312666
rect 563525 312632 563559 312640
rect 563525 312572 563559 312594
rect 563525 312560 563559 312572
rect 563525 312504 563559 312522
rect 563525 312488 563559 312504
rect 563525 312436 563559 312450
rect 563525 312416 563559 312436
rect 563525 312368 563559 312378
rect 563525 312344 563559 312368
rect 563525 312300 563559 312306
rect 563525 312272 563559 312300
rect 563525 312232 563559 312234
rect 563525 312200 563559 312232
rect 563525 312130 563559 312162
rect 563525 312128 563559 312130
rect 563525 312062 563559 312090
rect 563525 312056 563559 312062
rect 563525 311994 563559 312018
rect 563525 311984 563559 311994
rect 563525 311926 563559 311946
rect 563525 311912 563559 311926
rect 563525 311858 563559 311874
rect 563525 311840 563559 311858
rect 563525 311790 563559 311802
rect 563525 311768 563559 311790
rect 563525 311722 563559 311730
rect 563525 311696 563559 311722
rect 563783 312640 563817 312666
rect 563783 312632 563817 312640
rect 563783 312572 563817 312594
rect 563783 312560 563817 312572
rect 563783 312504 563817 312522
rect 563783 312488 563817 312504
rect 563783 312436 563817 312450
rect 563783 312416 563817 312436
rect 563783 312368 563817 312378
rect 563783 312344 563817 312368
rect 563783 312300 563817 312306
rect 563783 312272 563817 312300
rect 563783 312232 563817 312234
rect 563783 312200 563817 312232
rect 563783 312130 563817 312162
rect 563783 312128 563817 312130
rect 563783 312062 563817 312090
rect 563783 312056 563817 312062
rect 563783 311994 563817 312018
rect 563783 311984 563817 311994
rect 563783 311926 563817 311946
rect 563783 311912 563817 311926
rect 563783 311858 563817 311874
rect 563783 311840 563817 311858
rect 563783 311790 563817 311802
rect 563783 311768 563817 311790
rect 563783 311722 563817 311730
rect 563783 311696 563817 311722
rect 564041 312640 564075 312666
rect 564041 312632 564075 312640
rect 564041 312572 564075 312594
rect 564041 312560 564075 312572
rect 564041 312504 564075 312522
rect 564041 312488 564075 312504
rect 564041 312436 564075 312450
rect 564041 312416 564075 312436
rect 564041 312368 564075 312378
rect 564041 312344 564075 312368
rect 564041 312300 564075 312306
rect 564041 312272 564075 312300
rect 564041 312232 564075 312234
rect 564041 312200 564075 312232
rect 564041 312130 564075 312162
rect 564041 312128 564075 312130
rect 564041 312062 564075 312090
rect 564041 312056 564075 312062
rect 564041 311994 564075 312018
rect 564041 311984 564075 311994
rect 564041 311926 564075 311946
rect 564041 311912 564075 311926
rect 564041 311858 564075 311874
rect 564041 311840 564075 311858
rect 564041 311790 564075 311802
rect 564041 311768 564075 311790
rect 564041 311722 564075 311730
rect 564041 311696 564075 311722
rect 564299 312640 564333 312666
rect 564299 312632 564333 312640
rect 564299 312572 564333 312594
rect 564299 312560 564333 312572
rect 564299 312504 564333 312522
rect 564299 312488 564333 312504
rect 564299 312436 564333 312450
rect 564299 312416 564333 312436
rect 564299 312368 564333 312378
rect 564299 312344 564333 312368
rect 564299 312300 564333 312306
rect 564299 312272 564333 312300
rect 564299 312232 564333 312234
rect 564299 312200 564333 312232
rect 564299 312130 564333 312162
rect 564299 312128 564333 312130
rect 564299 312062 564333 312090
rect 564299 312056 564333 312062
rect 564299 311994 564333 312018
rect 564299 311984 564333 311994
rect 564299 311926 564333 311946
rect 564299 311912 564333 311926
rect 564299 311858 564333 311874
rect 564299 311840 564333 311858
rect 564299 311790 564333 311802
rect 564299 311768 564333 311790
rect 564299 311722 564333 311730
rect 564299 311696 564333 311722
rect 564557 312640 564591 312666
rect 564557 312632 564591 312640
rect 564557 312572 564591 312594
rect 564557 312560 564591 312572
rect 564557 312504 564591 312522
rect 564557 312488 564591 312504
rect 564557 312436 564591 312450
rect 564557 312416 564591 312436
rect 564557 312368 564591 312378
rect 564557 312344 564591 312368
rect 564557 312300 564591 312306
rect 564557 312272 564591 312300
rect 564557 312232 564591 312234
rect 564557 312200 564591 312232
rect 564557 312130 564591 312162
rect 564557 312128 564591 312130
rect 564557 312062 564591 312090
rect 564557 312056 564591 312062
rect 564557 311994 564591 312018
rect 564557 311984 564591 311994
rect 564557 311926 564591 311946
rect 564557 311912 564591 311926
rect 564557 311858 564591 311874
rect 564557 311840 564591 311858
rect 564557 311790 564591 311802
rect 564557 311768 564591 311790
rect 564557 311722 564591 311730
rect 564557 311696 564591 311722
rect 564815 312640 564849 312666
rect 564815 312632 564849 312640
rect 564815 312572 564849 312594
rect 564815 312560 564849 312572
rect 564815 312504 564849 312522
rect 564815 312488 564849 312504
rect 564815 312436 564849 312450
rect 564815 312416 564849 312436
rect 564815 312368 564849 312378
rect 564815 312344 564849 312368
rect 564815 312300 564849 312306
rect 564815 312272 564849 312300
rect 564815 312232 564849 312234
rect 564815 312200 564849 312232
rect 564815 312130 564849 312162
rect 564815 312128 564849 312130
rect 564815 312062 564849 312090
rect 564815 312056 564849 312062
rect 564815 311994 564849 312018
rect 564815 311984 564849 311994
rect 564815 311926 564849 311946
rect 564815 311912 564849 311926
rect 564815 311858 564849 311874
rect 564815 311840 564849 311858
rect 564815 311790 564849 311802
rect 564815 311768 564849 311790
rect 564815 311722 564849 311730
rect 564815 311696 564849 311722
rect 565073 312640 565107 312666
rect 565073 312632 565107 312640
rect 565073 312572 565107 312594
rect 565073 312560 565107 312572
rect 565073 312504 565107 312522
rect 565073 312488 565107 312504
rect 565073 312436 565107 312450
rect 565073 312416 565107 312436
rect 565073 312368 565107 312378
rect 565073 312344 565107 312368
rect 565073 312300 565107 312306
rect 565073 312272 565107 312300
rect 565073 312232 565107 312234
rect 565073 312200 565107 312232
rect 565073 312130 565107 312162
rect 565073 312128 565107 312130
rect 565073 312062 565107 312090
rect 565073 312056 565107 312062
rect 565073 311994 565107 312018
rect 565073 311984 565107 311994
rect 565073 311926 565107 311946
rect 565073 311912 565107 311926
rect 565073 311858 565107 311874
rect 565073 311840 565107 311858
rect 565073 311790 565107 311802
rect 565073 311768 565107 311790
rect 565073 311722 565107 311730
rect 565073 311696 565107 311722
rect 565331 312640 565365 312666
rect 565331 312632 565365 312640
rect 565331 312572 565365 312594
rect 565331 312560 565365 312572
rect 565331 312504 565365 312522
rect 565331 312488 565365 312504
rect 565331 312436 565365 312450
rect 565331 312416 565365 312436
rect 565331 312368 565365 312378
rect 565331 312344 565365 312368
rect 565331 312300 565365 312306
rect 565331 312272 565365 312300
rect 565331 312232 565365 312234
rect 565331 312200 565365 312232
rect 565331 312130 565365 312162
rect 565331 312128 565365 312130
rect 565331 312062 565365 312090
rect 565331 312056 565365 312062
rect 565331 311994 565365 312018
rect 565331 311984 565365 311994
rect 565331 311926 565365 311946
rect 565331 311912 565365 311926
rect 565331 311858 565365 311874
rect 565331 311840 565365 311858
rect 565331 311790 565365 311802
rect 565331 311768 565365 311790
rect 565331 311722 565365 311730
rect 565331 311696 565365 311722
rect 565589 312640 565623 312666
rect 565589 312632 565623 312640
rect 565589 312572 565623 312594
rect 565589 312560 565623 312572
rect 565589 312504 565623 312522
rect 565589 312488 565623 312504
rect 565589 312436 565623 312450
rect 565589 312416 565623 312436
rect 565589 312368 565623 312378
rect 565589 312344 565623 312368
rect 565589 312300 565623 312306
rect 565589 312272 565623 312300
rect 565589 312232 565623 312234
rect 565589 312200 565623 312232
rect 565589 312130 565623 312162
rect 565589 312128 565623 312130
rect 565589 312062 565623 312090
rect 565589 312056 565623 312062
rect 565589 311994 565623 312018
rect 565589 311984 565623 311994
rect 565589 311926 565623 311946
rect 565589 311912 565623 311926
rect 565589 311858 565623 311874
rect 565589 311840 565623 311858
rect 565589 311790 565623 311802
rect 565589 311768 565623 311790
rect 565589 311722 565623 311730
rect 565589 311696 565623 311722
rect 565869 311562 565975 311668
rect 575153 312710 575187 312736
rect 575153 312702 575187 312710
rect 575153 312642 575187 312664
rect 575153 312630 575187 312642
rect 575153 312574 575187 312592
rect 575153 312558 575187 312574
rect 575153 312506 575187 312520
rect 575153 312486 575187 312506
rect 575153 312438 575187 312448
rect 575153 312414 575187 312438
rect 575153 312370 575187 312376
rect 575153 312342 575187 312370
rect 575153 312302 575187 312304
rect 575153 312270 575187 312302
rect 575153 312200 575187 312232
rect 575153 312198 575187 312200
rect 575153 312132 575187 312160
rect 575153 312126 575187 312132
rect 575153 312064 575187 312088
rect 575153 312054 575187 312064
rect 575153 311996 575187 312016
rect 575153 311982 575187 311996
rect 575153 311928 575187 311944
rect 575153 311910 575187 311928
rect 575153 311860 575187 311872
rect 575153 311838 575187 311860
rect 575153 311792 575187 311800
rect 575153 311766 575187 311792
rect 575411 312710 575445 312736
rect 575411 312702 575445 312710
rect 575411 312642 575445 312664
rect 575411 312630 575445 312642
rect 575411 312574 575445 312592
rect 575411 312558 575445 312574
rect 575411 312506 575445 312520
rect 575411 312486 575445 312506
rect 575411 312438 575445 312448
rect 575411 312414 575445 312438
rect 575411 312370 575445 312376
rect 575411 312342 575445 312370
rect 575411 312302 575445 312304
rect 575411 312270 575445 312302
rect 575411 312200 575445 312232
rect 575411 312198 575445 312200
rect 575411 312132 575445 312160
rect 575411 312126 575445 312132
rect 575411 312064 575445 312088
rect 575411 312054 575445 312064
rect 575411 311996 575445 312016
rect 575411 311982 575445 311996
rect 575411 311928 575445 311944
rect 575411 311910 575445 311928
rect 575411 311860 575445 311872
rect 575411 311838 575445 311860
rect 575411 311792 575445 311800
rect 575411 311766 575445 311792
rect 575669 312710 575703 312736
rect 575669 312702 575703 312710
rect 575669 312642 575703 312664
rect 575669 312630 575703 312642
rect 575669 312574 575703 312592
rect 575669 312558 575703 312574
rect 575669 312506 575703 312520
rect 575669 312486 575703 312506
rect 575669 312438 575703 312448
rect 575669 312414 575703 312438
rect 575669 312370 575703 312376
rect 575669 312342 575703 312370
rect 575669 312302 575703 312304
rect 575669 312270 575703 312302
rect 575669 312200 575703 312232
rect 575669 312198 575703 312200
rect 575669 312132 575703 312160
rect 575669 312126 575703 312132
rect 575669 312064 575703 312088
rect 575669 312054 575703 312064
rect 575669 311996 575703 312016
rect 575669 311982 575703 311996
rect 575669 311928 575703 311944
rect 575669 311910 575703 311928
rect 575669 311860 575703 311872
rect 575669 311838 575703 311860
rect 575669 311792 575703 311800
rect 575669 311766 575703 311792
rect 575927 312710 575961 312736
rect 575927 312702 575961 312710
rect 575927 312642 575961 312664
rect 575927 312630 575961 312642
rect 575927 312574 575961 312592
rect 575927 312558 575961 312574
rect 575927 312506 575961 312520
rect 575927 312486 575961 312506
rect 575927 312438 575961 312448
rect 575927 312414 575961 312438
rect 575927 312370 575961 312376
rect 575927 312342 575961 312370
rect 575927 312302 575961 312304
rect 575927 312270 575961 312302
rect 575927 312200 575961 312232
rect 575927 312198 575961 312200
rect 575927 312132 575961 312160
rect 575927 312126 575961 312132
rect 575927 312064 575961 312088
rect 575927 312054 575961 312064
rect 575927 311996 575961 312016
rect 575927 311982 575961 311996
rect 575927 311928 575961 311944
rect 575927 311910 575961 311928
rect 575927 311860 575961 311872
rect 575927 311838 575961 311860
rect 575927 311792 575961 311800
rect 575927 311766 575961 311792
rect 576185 312710 576219 312736
rect 576185 312702 576219 312710
rect 576185 312642 576219 312664
rect 576185 312630 576219 312642
rect 576185 312574 576219 312592
rect 576185 312558 576219 312574
rect 576185 312506 576219 312520
rect 576185 312486 576219 312506
rect 576185 312438 576219 312448
rect 576185 312414 576219 312438
rect 576185 312370 576219 312376
rect 576185 312342 576219 312370
rect 576185 312302 576219 312304
rect 576185 312270 576219 312302
rect 576185 312200 576219 312232
rect 576185 312198 576219 312200
rect 576185 312132 576219 312160
rect 576185 312126 576219 312132
rect 576185 312064 576219 312088
rect 576185 312054 576219 312064
rect 576185 311996 576219 312016
rect 576185 311982 576219 311996
rect 576185 311928 576219 311944
rect 576185 311910 576219 311928
rect 576185 311860 576219 311872
rect 576185 311838 576219 311860
rect 576185 311792 576219 311800
rect 576185 311766 576219 311792
rect 576443 312710 576477 312736
rect 576443 312702 576477 312710
rect 576443 312642 576477 312664
rect 576443 312630 576477 312642
rect 576443 312574 576477 312592
rect 576443 312558 576477 312574
rect 576443 312506 576477 312520
rect 576443 312486 576477 312506
rect 576443 312438 576477 312448
rect 576443 312414 576477 312438
rect 576443 312370 576477 312376
rect 576443 312342 576477 312370
rect 576443 312302 576477 312304
rect 576443 312270 576477 312302
rect 576443 312200 576477 312232
rect 576443 312198 576477 312200
rect 576443 312132 576477 312160
rect 576443 312126 576477 312132
rect 576443 312064 576477 312088
rect 576443 312054 576477 312064
rect 576443 311996 576477 312016
rect 576443 311982 576477 311996
rect 576443 311928 576477 311944
rect 576443 311910 576477 311928
rect 576443 311860 576477 311872
rect 576443 311838 576477 311860
rect 576443 311792 576477 311800
rect 576443 311766 576477 311792
rect 576701 312710 576735 312736
rect 576701 312702 576735 312710
rect 576701 312642 576735 312664
rect 576701 312630 576735 312642
rect 576701 312574 576735 312592
rect 576701 312558 576735 312574
rect 576701 312506 576735 312520
rect 576701 312486 576735 312506
rect 576701 312438 576735 312448
rect 576701 312414 576735 312438
rect 576701 312370 576735 312376
rect 576701 312342 576735 312370
rect 576701 312302 576735 312304
rect 576701 312270 576735 312302
rect 576701 312200 576735 312232
rect 576701 312198 576735 312200
rect 576701 312132 576735 312160
rect 576701 312126 576735 312132
rect 576701 312064 576735 312088
rect 576701 312054 576735 312064
rect 576701 311996 576735 312016
rect 576701 311982 576735 311996
rect 576701 311928 576735 311944
rect 576701 311910 576735 311928
rect 576701 311860 576735 311872
rect 576701 311838 576735 311860
rect 576701 311792 576735 311800
rect 576701 311766 576735 311792
rect 576959 312710 576993 312736
rect 576959 312702 576993 312710
rect 576959 312642 576993 312664
rect 576959 312630 576993 312642
rect 576959 312574 576993 312592
rect 576959 312558 576993 312574
rect 576959 312506 576993 312520
rect 576959 312486 576993 312506
rect 576959 312438 576993 312448
rect 576959 312414 576993 312438
rect 576959 312370 576993 312376
rect 576959 312342 576993 312370
rect 576959 312302 576993 312304
rect 576959 312270 576993 312302
rect 576959 312200 576993 312232
rect 576959 312198 576993 312200
rect 576959 312132 576993 312160
rect 576959 312126 576993 312132
rect 576959 312064 576993 312088
rect 576959 312054 576993 312064
rect 576959 311996 576993 312016
rect 576959 311982 576993 311996
rect 576959 311928 576993 311944
rect 576959 311910 576993 311928
rect 576959 311860 576993 311872
rect 576959 311838 576993 311860
rect 576959 311792 576993 311800
rect 576959 311766 576993 311792
rect 577217 312710 577251 312736
rect 577217 312702 577251 312710
rect 577217 312642 577251 312664
rect 577217 312630 577251 312642
rect 577217 312574 577251 312592
rect 577217 312558 577251 312574
rect 577217 312506 577251 312520
rect 577217 312486 577251 312506
rect 577217 312438 577251 312448
rect 577217 312414 577251 312438
rect 577217 312370 577251 312376
rect 577217 312342 577251 312370
rect 577217 312302 577251 312304
rect 577217 312270 577251 312302
rect 577217 312200 577251 312232
rect 577217 312198 577251 312200
rect 577217 312132 577251 312160
rect 577217 312126 577251 312132
rect 577217 312064 577251 312088
rect 577217 312054 577251 312064
rect 577217 311996 577251 312016
rect 577217 311982 577251 311996
rect 577217 311928 577251 311944
rect 577217 311910 577251 311928
rect 577217 311860 577251 311872
rect 577217 311838 577251 311860
rect 577217 311792 577251 311800
rect 577217 311766 577251 311792
rect 577475 312710 577509 312736
rect 577475 312702 577509 312710
rect 577475 312642 577509 312664
rect 577475 312630 577509 312642
rect 577475 312574 577509 312592
rect 577475 312558 577509 312574
rect 577475 312506 577509 312520
rect 577475 312486 577509 312506
rect 577475 312438 577509 312448
rect 577475 312414 577509 312438
rect 577475 312370 577509 312376
rect 577475 312342 577509 312370
rect 577475 312302 577509 312304
rect 577475 312270 577509 312302
rect 577475 312200 577509 312232
rect 577475 312198 577509 312200
rect 577475 312132 577509 312160
rect 577475 312126 577509 312132
rect 577475 312064 577509 312088
rect 577475 312054 577509 312064
rect 577475 311996 577509 312016
rect 577475 311982 577509 311996
rect 577475 311928 577509 311944
rect 577475 311910 577509 311928
rect 577475 311860 577509 311872
rect 577475 311838 577509 311860
rect 577475 311792 577509 311800
rect 577475 311766 577509 311792
rect 577733 312710 577767 312736
rect 577733 312702 577767 312710
rect 577733 312642 577767 312664
rect 577733 312630 577767 312642
rect 577733 312574 577767 312592
rect 577733 312558 577767 312574
rect 577733 312506 577767 312520
rect 577733 312486 577767 312506
rect 577733 312438 577767 312448
rect 577733 312414 577767 312438
rect 577733 312370 577767 312376
rect 577733 312342 577767 312370
rect 577733 312302 577767 312304
rect 577733 312270 577767 312302
rect 577733 312200 577767 312232
rect 577733 312198 577767 312200
rect 577733 312132 577767 312160
rect 577733 312126 577767 312132
rect 577733 312064 577767 312088
rect 577733 312054 577767 312064
rect 577733 311996 577767 312016
rect 577733 311982 577767 311996
rect 577733 311928 577767 311944
rect 577733 311910 577767 311928
rect 577733 311860 577767 311872
rect 577733 311838 577767 311860
rect 577733 311792 577767 311800
rect 577733 311766 577767 311792
rect 577991 312710 578025 312736
rect 577991 312702 578025 312710
rect 577991 312642 578025 312664
rect 577991 312630 578025 312642
rect 577991 312574 578025 312592
rect 577991 312558 578025 312574
rect 577991 312506 578025 312520
rect 577991 312486 578025 312506
rect 577991 312438 578025 312448
rect 577991 312414 578025 312438
rect 577991 312370 578025 312376
rect 577991 312342 578025 312370
rect 577991 312302 578025 312304
rect 577991 312270 578025 312302
rect 577991 312200 578025 312232
rect 577991 312198 578025 312200
rect 577991 312132 578025 312160
rect 577991 312126 578025 312132
rect 577991 312064 578025 312088
rect 577991 312054 578025 312064
rect 577991 311996 578025 312016
rect 577991 311982 578025 311996
rect 577991 311928 578025 311944
rect 577991 311910 578025 311928
rect 577991 311860 578025 311872
rect 577991 311838 578025 311860
rect 577991 311792 578025 311800
rect 577991 311766 578025 311792
rect 578249 312710 578283 312736
rect 578249 312702 578283 312710
rect 578249 312642 578283 312664
rect 578249 312630 578283 312642
rect 578249 312574 578283 312592
rect 578249 312558 578283 312574
rect 578249 312506 578283 312520
rect 578249 312486 578283 312506
rect 578249 312438 578283 312448
rect 578249 312414 578283 312438
rect 578249 312370 578283 312376
rect 578249 312342 578283 312370
rect 578249 312302 578283 312304
rect 578249 312270 578283 312302
rect 578249 312200 578283 312232
rect 578249 312198 578283 312200
rect 578249 312132 578283 312160
rect 578249 312126 578283 312132
rect 578249 312064 578283 312088
rect 578249 312054 578283 312064
rect 578249 311996 578283 312016
rect 578249 311982 578283 311996
rect 578249 311928 578283 311944
rect 578249 311910 578283 311928
rect 578249 311860 578283 311872
rect 578249 311838 578283 311860
rect 578249 311792 578283 311800
rect 578249 311766 578283 311792
rect 578507 312710 578541 312736
rect 578507 312702 578541 312710
rect 578507 312642 578541 312664
rect 578507 312630 578541 312642
rect 578507 312574 578541 312592
rect 578507 312558 578541 312574
rect 578507 312506 578541 312520
rect 578507 312486 578541 312506
rect 578507 312438 578541 312448
rect 578507 312414 578541 312438
rect 578507 312370 578541 312376
rect 578507 312342 578541 312370
rect 578507 312302 578541 312304
rect 578507 312270 578541 312302
rect 578507 312200 578541 312232
rect 578507 312198 578541 312200
rect 578507 312132 578541 312160
rect 578507 312126 578541 312132
rect 578507 312064 578541 312088
rect 578507 312054 578541 312064
rect 578507 311996 578541 312016
rect 578507 311982 578541 311996
rect 578507 311928 578541 311944
rect 578507 311910 578541 311928
rect 578507 311860 578541 311872
rect 578507 311838 578541 311860
rect 578507 311792 578541 311800
rect 578507 311766 578541 311792
rect 578765 312710 578799 312736
rect 578765 312702 578799 312710
rect 578765 312642 578799 312664
rect 578765 312630 578799 312642
rect 578765 312574 578799 312592
rect 578765 312558 578799 312574
rect 578765 312506 578799 312520
rect 578765 312486 578799 312506
rect 578765 312438 578799 312448
rect 578765 312414 578799 312438
rect 578765 312370 578799 312376
rect 578765 312342 578799 312370
rect 578765 312302 578799 312304
rect 578765 312270 578799 312302
rect 578765 312200 578799 312232
rect 578765 312198 578799 312200
rect 578765 312132 578799 312160
rect 578765 312126 578799 312132
rect 578765 312064 578799 312088
rect 578765 312054 578799 312064
rect 578765 311996 578799 312016
rect 578765 311982 578799 311996
rect 578765 311928 578799 311944
rect 578765 311910 578799 311928
rect 578765 311860 578799 311872
rect 578765 311838 578799 311860
rect 578765 311792 578799 311800
rect 578765 311766 578799 311792
rect 579023 312710 579057 312736
rect 579023 312702 579057 312710
rect 579023 312642 579057 312664
rect 579023 312630 579057 312642
rect 579023 312574 579057 312592
rect 579023 312558 579057 312574
rect 579023 312506 579057 312520
rect 579023 312486 579057 312506
rect 579023 312438 579057 312448
rect 579023 312414 579057 312438
rect 579023 312370 579057 312376
rect 579023 312342 579057 312370
rect 579023 312302 579057 312304
rect 579023 312270 579057 312302
rect 579023 312200 579057 312232
rect 579023 312198 579057 312200
rect 579023 312132 579057 312160
rect 579023 312126 579057 312132
rect 579023 312064 579057 312088
rect 579023 312054 579057 312064
rect 579023 311996 579057 312016
rect 579023 311982 579057 311996
rect 579023 311928 579057 311944
rect 579023 311910 579057 311928
rect 579023 311860 579057 311872
rect 579023 311838 579057 311860
rect 579023 311792 579057 311800
rect 579023 311766 579057 311792
rect 579281 312710 579315 312736
rect 579281 312702 579315 312710
rect 579281 312642 579315 312664
rect 579281 312630 579315 312642
rect 579281 312574 579315 312592
rect 579281 312558 579315 312574
rect 579281 312506 579315 312520
rect 579281 312486 579315 312506
rect 579281 312438 579315 312448
rect 579281 312414 579315 312438
rect 579281 312370 579315 312376
rect 579281 312342 579315 312370
rect 579281 312302 579315 312304
rect 579281 312270 579315 312302
rect 579281 312200 579315 312232
rect 579281 312198 579315 312200
rect 579281 312132 579315 312160
rect 579281 312126 579315 312132
rect 579281 312064 579315 312088
rect 579281 312054 579315 312064
rect 579281 311996 579315 312016
rect 579281 311982 579315 311996
rect 579281 311928 579315 311944
rect 579281 311910 579315 311928
rect 579281 311860 579315 311872
rect 579281 311838 579315 311860
rect 579281 311792 579315 311800
rect 579281 311766 579315 311792
rect 579539 312710 579573 312736
rect 579539 312702 579573 312710
rect 579539 312642 579573 312664
rect 579539 312630 579573 312642
rect 579539 312574 579573 312592
rect 579539 312558 579573 312574
rect 579539 312506 579573 312520
rect 579539 312486 579573 312506
rect 579539 312438 579573 312448
rect 579539 312414 579573 312438
rect 579539 312370 579573 312376
rect 579539 312342 579573 312370
rect 579539 312302 579573 312304
rect 579539 312270 579573 312302
rect 579539 312200 579573 312232
rect 579539 312198 579573 312200
rect 579539 312132 579573 312160
rect 579539 312126 579573 312132
rect 579539 312064 579573 312088
rect 579539 312054 579573 312064
rect 579539 311996 579573 312016
rect 579539 311982 579573 311996
rect 579539 311928 579573 311944
rect 579539 311910 579573 311928
rect 579539 311860 579573 311872
rect 579539 311838 579573 311860
rect 579539 311792 579573 311800
rect 579539 311766 579573 311792
rect 579797 312710 579831 312736
rect 579797 312702 579831 312710
rect 579797 312642 579831 312664
rect 579797 312630 579831 312642
rect 579797 312574 579831 312592
rect 579797 312558 579831 312574
rect 579797 312506 579831 312520
rect 579797 312486 579831 312506
rect 579797 312438 579831 312448
rect 579797 312414 579831 312438
rect 579797 312370 579831 312376
rect 579797 312342 579831 312370
rect 579797 312302 579831 312304
rect 579797 312270 579831 312302
rect 579797 312200 579831 312232
rect 579797 312198 579831 312200
rect 579797 312132 579831 312160
rect 579797 312126 579831 312132
rect 579797 312064 579831 312088
rect 579797 312054 579831 312064
rect 579797 311996 579831 312016
rect 579797 311982 579831 311996
rect 579797 311928 579831 311944
rect 579797 311910 579831 311928
rect 579797 311860 579831 311872
rect 579797 311838 579831 311860
rect 579797 311792 579831 311800
rect 579797 311766 579831 311792
rect 580055 312710 580089 312736
rect 580055 312702 580089 312710
rect 580055 312642 580089 312664
rect 580055 312630 580089 312642
rect 580055 312574 580089 312592
rect 580055 312558 580089 312574
rect 580055 312506 580089 312520
rect 580055 312486 580089 312506
rect 580055 312438 580089 312448
rect 580055 312414 580089 312438
rect 580055 312370 580089 312376
rect 580055 312342 580089 312370
rect 580055 312302 580089 312304
rect 580055 312270 580089 312302
rect 580055 312200 580089 312232
rect 580055 312198 580089 312200
rect 580055 312132 580089 312160
rect 580055 312126 580089 312132
rect 580055 312064 580089 312088
rect 580055 312054 580089 312064
rect 580055 311996 580089 312016
rect 580055 311982 580089 311996
rect 580055 311928 580089 311944
rect 580055 311910 580089 311928
rect 580055 311860 580089 311872
rect 580055 311838 580089 311860
rect 580055 311792 580089 311800
rect 580055 311766 580089 311792
rect 580313 312710 580347 312736
rect 580313 312702 580347 312710
rect 580313 312642 580347 312664
rect 580313 312630 580347 312642
rect 580313 312574 580347 312592
rect 580313 312558 580347 312574
rect 580313 312506 580347 312520
rect 580313 312486 580347 312506
rect 580313 312438 580347 312448
rect 580313 312414 580347 312438
rect 580313 312370 580347 312376
rect 580313 312342 580347 312370
rect 580313 312302 580347 312304
rect 580313 312270 580347 312302
rect 580313 312200 580347 312232
rect 580313 312198 580347 312200
rect 580313 312132 580347 312160
rect 580313 312126 580347 312132
rect 580313 312064 580347 312088
rect 580313 312054 580347 312064
rect 580313 311996 580347 312016
rect 580313 311982 580347 311996
rect 580313 311928 580347 311944
rect 580313 311910 580347 311928
rect 580313 311860 580347 311872
rect 580313 311838 580347 311860
rect 580313 311792 580347 311800
rect 580313 311766 580347 311792
rect 580506 311594 580540 311628
rect 574899 311452 574933 311486
rect 575177 311234 575211 311268
rect 575377 311234 575411 311268
rect 575577 311234 575611 311268
rect 575777 311234 575811 311268
rect 575977 311234 576011 311268
rect 576177 311234 576211 311268
rect 576377 311234 576411 311268
rect 576577 311234 576611 311268
rect 576777 311234 576811 311268
rect 576977 311234 577011 311268
rect 577177 311234 577211 311268
rect 577377 311234 577411 311268
rect 577577 311234 577611 311268
rect 577777 311234 577811 311268
rect 577977 311234 578011 311268
rect 578177 311234 578211 311268
rect 578377 311234 578411 311268
rect 578577 311234 578611 311268
rect 578777 311234 578811 311268
rect 578977 311234 579011 311268
rect 579177 311234 579211 311268
rect 579377 311234 579411 311268
rect 579577 311234 579611 311268
rect 579777 311234 579811 311268
rect 579977 311234 580011 311268
rect 580177 311234 580211 311268
rect 560617 311164 560651 311198
rect 560817 311164 560851 311198
rect 561017 311164 561051 311198
rect 561217 311164 561251 311198
rect 561417 311164 561451 311198
rect 561617 311164 561651 311198
rect 561817 311164 561851 311198
rect 562017 311164 562051 311198
rect 562217 311164 562251 311198
rect 562417 311164 562451 311198
rect 562617 311164 562651 311198
rect 562817 311164 562851 311198
rect 563017 311164 563051 311198
rect 563217 311164 563251 311198
rect 563417 311164 563451 311198
rect 563617 311164 563651 311198
rect 563817 311164 563851 311198
rect 564017 311164 564051 311198
rect 564217 311164 564251 311198
rect 564417 311164 564451 311198
rect 564617 311164 564651 311198
rect 564817 311164 564851 311198
rect 565017 311164 565051 311198
rect 565217 311164 565251 311198
rect 565417 311164 565451 311198
<< metal1 >>
rect 573598 494891 573810 494897
rect 565710 494771 573810 494891
rect 565710 493889 565830 494771
rect 566190 494317 566432 494319
rect 566190 494137 566221 494317
rect 566401 494137 566432 494317
rect 566190 494135 566432 494137
rect 560664 493846 565978 493889
rect 560664 493812 560863 493846
rect 560897 493812 561063 493846
rect 561097 493812 561263 493846
rect 561297 493812 561463 493846
rect 561497 493812 561663 493846
rect 561697 493812 561863 493846
rect 561897 493812 562063 493846
rect 562097 493812 562263 493846
rect 562297 493812 562463 493846
rect 562497 493812 562663 493846
rect 562697 493812 562863 493846
rect 562897 493812 563063 493846
rect 563097 493812 563263 493846
rect 563297 493812 563463 493846
rect 563497 493812 563663 493846
rect 563697 493812 563863 493846
rect 563897 493812 564063 493846
rect 564097 493812 564263 493846
rect 564297 493812 564463 493846
rect 564497 493812 564663 493846
rect 564697 493812 564863 493846
rect 564897 493812 565063 493846
rect 565097 493812 565263 493846
rect 565297 493812 565463 493846
rect 565497 493812 565663 493846
rect 565697 493812 565978 493846
rect 560664 493769 565978 493812
rect 560669 493434 560715 493449
rect 560669 493400 560675 493434
rect 560709 493400 560715 493434
rect 560669 493362 560715 493400
rect 560669 493328 560675 493362
rect 560709 493328 560715 493362
rect 560669 493290 560715 493328
rect 560669 493256 560675 493290
rect 560709 493256 560715 493290
rect 560669 493218 560715 493256
rect 560669 493184 560675 493218
rect 560709 493184 560715 493218
rect 560669 493146 560715 493184
rect 560669 493112 560675 493146
rect 560709 493112 560715 493146
rect 560669 493074 560715 493112
rect 560669 493040 560675 493074
rect 560709 493040 560715 493074
rect 560669 493002 560715 493040
rect 560669 492968 560675 493002
rect 560709 492968 560715 493002
rect 560669 492930 560715 492968
rect 560669 492896 560675 492930
rect 560709 492896 560715 492930
rect 560669 492858 560715 492896
rect 560669 492824 560675 492858
rect 560709 492824 560715 492858
rect 560669 492786 560715 492824
rect 560669 492752 560675 492786
rect 560709 492752 560715 492786
rect 560669 492714 560715 492752
rect 560669 492680 560675 492714
rect 560709 492680 560715 492714
rect 560669 492642 560715 492680
rect 560669 492608 560675 492642
rect 560709 492608 560715 492642
rect 560669 492570 560715 492608
rect 559806 492557 560124 492563
rect 559802 492529 560462 492557
rect 559802 492349 559831 492529
rect 560011 492521 560462 492529
rect 560669 492536 560675 492570
rect 560709 492536 560715 492570
rect 560011 492469 560500 492521
rect 560011 492363 560367 492469
rect 560473 492363 560500 492469
rect 560669 492498 560715 492536
rect 560669 492464 560675 492498
rect 560709 492464 560715 492498
rect 560669 492449 560715 492464
rect 560927 493434 560973 493449
rect 560927 493400 560933 493434
rect 560967 493400 560973 493434
rect 560927 493362 560973 493400
rect 560927 493328 560933 493362
rect 560967 493328 560973 493362
rect 560927 493290 560973 493328
rect 560927 493256 560933 493290
rect 560967 493256 560973 493290
rect 560927 493218 560973 493256
rect 560927 493184 560933 493218
rect 560967 493184 560973 493218
rect 560927 493146 560973 493184
rect 560927 493112 560933 493146
rect 560967 493112 560973 493146
rect 560927 493074 560973 493112
rect 560927 493040 560933 493074
rect 560967 493040 560973 493074
rect 560927 493002 560973 493040
rect 560927 492968 560933 493002
rect 560967 492968 560973 493002
rect 560927 492930 560973 492968
rect 560927 492896 560933 492930
rect 560967 492896 560973 492930
rect 560927 492858 560973 492896
rect 560927 492824 560933 492858
rect 560967 492824 560973 492858
rect 560927 492786 560973 492824
rect 560927 492752 560933 492786
rect 560967 492752 560973 492786
rect 560927 492714 560973 492752
rect 560927 492680 560933 492714
rect 560967 492680 560973 492714
rect 560927 492642 560973 492680
rect 560927 492608 560933 492642
rect 560967 492608 560973 492642
rect 560927 492570 560973 492608
rect 560927 492536 560933 492570
rect 560967 492536 560973 492570
rect 560927 492498 560973 492536
rect 560927 492464 560933 492498
rect 560967 492464 560973 492498
rect 560927 492449 560973 492464
rect 561185 493434 561231 493449
rect 561185 493400 561191 493434
rect 561225 493400 561231 493434
rect 561185 493362 561231 493400
rect 561185 493328 561191 493362
rect 561225 493328 561231 493362
rect 561185 493290 561231 493328
rect 561185 493256 561191 493290
rect 561225 493256 561231 493290
rect 561185 493218 561231 493256
rect 561185 493184 561191 493218
rect 561225 493184 561231 493218
rect 561185 493146 561231 493184
rect 561185 493112 561191 493146
rect 561225 493112 561231 493146
rect 561185 493074 561231 493112
rect 561185 493040 561191 493074
rect 561225 493040 561231 493074
rect 561185 493002 561231 493040
rect 561185 492968 561191 493002
rect 561225 492968 561231 493002
rect 561185 492930 561231 492968
rect 561185 492896 561191 492930
rect 561225 492896 561231 492930
rect 561185 492858 561231 492896
rect 561185 492824 561191 492858
rect 561225 492824 561231 492858
rect 561185 492786 561231 492824
rect 561185 492752 561191 492786
rect 561225 492752 561231 492786
rect 561185 492714 561231 492752
rect 561185 492680 561191 492714
rect 561225 492680 561231 492714
rect 561185 492642 561231 492680
rect 561185 492608 561191 492642
rect 561225 492608 561231 492642
rect 561185 492570 561231 492608
rect 561185 492536 561191 492570
rect 561225 492536 561231 492570
rect 561185 492498 561231 492536
rect 561185 492464 561191 492498
rect 561225 492464 561231 492498
rect 561185 492449 561231 492464
rect 561443 493434 561489 493449
rect 561443 493400 561449 493434
rect 561483 493400 561489 493434
rect 561443 493362 561489 493400
rect 561443 493328 561449 493362
rect 561483 493328 561489 493362
rect 561443 493290 561489 493328
rect 561443 493256 561449 493290
rect 561483 493256 561489 493290
rect 561443 493218 561489 493256
rect 561443 493184 561449 493218
rect 561483 493184 561489 493218
rect 561443 493146 561489 493184
rect 561443 493112 561449 493146
rect 561483 493112 561489 493146
rect 561443 493074 561489 493112
rect 561443 493040 561449 493074
rect 561483 493040 561489 493074
rect 561443 493002 561489 493040
rect 561443 492968 561449 493002
rect 561483 492968 561489 493002
rect 561443 492930 561489 492968
rect 561443 492896 561449 492930
rect 561483 492896 561489 492930
rect 561443 492858 561489 492896
rect 561443 492824 561449 492858
rect 561483 492824 561489 492858
rect 561443 492786 561489 492824
rect 561443 492752 561449 492786
rect 561483 492752 561489 492786
rect 561443 492714 561489 492752
rect 561443 492680 561449 492714
rect 561483 492680 561489 492714
rect 561443 492642 561489 492680
rect 561443 492608 561449 492642
rect 561483 492608 561489 492642
rect 561443 492570 561489 492608
rect 561443 492536 561449 492570
rect 561483 492536 561489 492570
rect 561443 492498 561489 492536
rect 561443 492464 561449 492498
rect 561483 492464 561489 492498
rect 561443 492449 561489 492464
rect 561701 493434 561747 493449
rect 561701 493400 561707 493434
rect 561741 493400 561747 493434
rect 561701 493362 561747 493400
rect 561701 493328 561707 493362
rect 561741 493328 561747 493362
rect 561701 493290 561747 493328
rect 561701 493256 561707 493290
rect 561741 493256 561747 493290
rect 561701 493218 561747 493256
rect 561701 493184 561707 493218
rect 561741 493184 561747 493218
rect 561701 493146 561747 493184
rect 561701 493112 561707 493146
rect 561741 493112 561747 493146
rect 561701 493074 561747 493112
rect 561701 493040 561707 493074
rect 561741 493040 561747 493074
rect 561701 493002 561747 493040
rect 561701 492968 561707 493002
rect 561741 492968 561747 493002
rect 561701 492930 561747 492968
rect 561701 492896 561707 492930
rect 561741 492896 561747 492930
rect 561701 492858 561747 492896
rect 561701 492824 561707 492858
rect 561741 492824 561747 492858
rect 561701 492786 561747 492824
rect 561701 492752 561707 492786
rect 561741 492752 561747 492786
rect 561701 492714 561747 492752
rect 561701 492680 561707 492714
rect 561741 492680 561747 492714
rect 561701 492642 561747 492680
rect 561701 492608 561707 492642
rect 561741 492608 561747 492642
rect 561701 492570 561747 492608
rect 561701 492536 561707 492570
rect 561741 492536 561747 492570
rect 561701 492498 561747 492536
rect 561701 492464 561707 492498
rect 561741 492464 561747 492498
rect 561701 492449 561747 492464
rect 561959 493434 562005 493449
rect 561959 493400 561965 493434
rect 561999 493400 562005 493434
rect 561959 493362 562005 493400
rect 561959 493328 561965 493362
rect 561999 493328 562005 493362
rect 561959 493290 562005 493328
rect 561959 493256 561965 493290
rect 561999 493256 562005 493290
rect 561959 493218 562005 493256
rect 561959 493184 561965 493218
rect 561999 493184 562005 493218
rect 561959 493146 562005 493184
rect 561959 493112 561965 493146
rect 561999 493112 562005 493146
rect 561959 493074 562005 493112
rect 561959 493040 561965 493074
rect 561999 493040 562005 493074
rect 561959 493002 562005 493040
rect 561959 492968 561965 493002
rect 561999 492968 562005 493002
rect 561959 492930 562005 492968
rect 561959 492896 561965 492930
rect 561999 492896 562005 492930
rect 561959 492858 562005 492896
rect 561959 492824 561965 492858
rect 561999 492824 562005 492858
rect 561959 492786 562005 492824
rect 561959 492752 561965 492786
rect 561999 492752 562005 492786
rect 561959 492714 562005 492752
rect 561959 492680 561965 492714
rect 561999 492680 562005 492714
rect 561959 492642 562005 492680
rect 561959 492608 561965 492642
rect 561999 492608 562005 492642
rect 561959 492570 562005 492608
rect 561959 492536 561965 492570
rect 561999 492536 562005 492570
rect 561959 492498 562005 492536
rect 561959 492464 561965 492498
rect 561999 492464 562005 492498
rect 561959 492449 562005 492464
rect 562217 493434 562263 493449
rect 562217 493400 562223 493434
rect 562257 493400 562263 493434
rect 562217 493362 562263 493400
rect 562217 493328 562223 493362
rect 562257 493328 562263 493362
rect 562217 493290 562263 493328
rect 562217 493256 562223 493290
rect 562257 493256 562263 493290
rect 562217 493218 562263 493256
rect 562217 493184 562223 493218
rect 562257 493184 562263 493218
rect 562217 493146 562263 493184
rect 562217 493112 562223 493146
rect 562257 493112 562263 493146
rect 562217 493074 562263 493112
rect 562217 493040 562223 493074
rect 562257 493040 562263 493074
rect 562217 493002 562263 493040
rect 562217 492968 562223 493002
rect 562257 492968 562263 493002
rect 562217 492930 562263 492968
rect 562217 492896 562223 492930
rect 562257 492896 562263 492930
rect 562217 492858 562263 492896
rect 562217 492824 562223 492858
rect 562257 492824 562263 492858
rect 562217 492786 562263 492824
rect 562217 492752 562223 492786
rect 562257 492752 562263 492786
rect 562217 492714 562263 492752
rect 562217 492680 562223 492714
rect 562257 492680 562263 492714
rect 562217 492642 562263 492680
rect 562217 492608 562223 492642
rect 562257 492608 562263 492642
rect 562217 492570 562263 492608
rect 562217 492536 562223 492570
rect 562257 492536 562263 492570
rect 562217 492498 562263 492536
rect 562217 492464 562223 492498
rect 562257 492464 562263 492498
rect 562217 492449 562263 492464
rect 562475 493434 562521 493449
rect 562475 493400 562481 493434
rect 562515 493400 562521 493434
rect 562475 493362 562521 493400
rect 562475 493328 562481 493362
rect 562515 493328 562521 493362
rect 562475 493290 562521 493328
rect 562475 493256 562481 493290
rect 562515 493256 562521 493290
rect 562475 493218 562521 493256
rect 562475 493184 562481 493218
rect 562515 493184 562521 493218
rect 562475 493146 562521 493184
rect 562475 493112 562481 493146
rect 562515 493112 562521 493146
rect 562475 493074 562521 493112
rect 562475 493040 562481 493074
rect 562515 493040 562521 493074
rect 562475 493002 562521 493040
rect 562475 492968 562481 493002
rect 562515 492968 562521 493002
rect 562475 492930 562521 492968
rect 562475 492896 562481 492930
rect 562515 492896 562521 492930
rect 562475 492858 562521 492896
rect 562475 492824 562481 492858
rect 562515 492824 562521 492858
rect 562475 492786 562521 492824
rect 562475 492752 562481 492786
rect 562515 492752 562521 492786
rect 562475 492714 562521 492752
rect 562475 492680 562481 492714
rect 562515 492680 562521 492714
rect 562475 492642 562521 492680
rect 562475 492608 562481 492642
rect 562515 492608 562521 492642
rect 562475 492570 562521 492608
rect 562475 492536 562481 492570
rect 562515 492536 562521 492570
rect 562475 492498 562521 492536
rect 562475 492464 562481 492498
rect 562515 492464 562521 492498
rect 562475 492449 562521 492464
rect 562733 493434 562779 493449
rect 562733 493400 562739 493434
rect 562773 493400 562779 493434
rect 562733 493362 562779 493400
rect 562733 493328 562739 493362
rect 562773 493328 562779 493362
rect 562733 493290 562779 493328
rect 562733 493256 562739 493290
rect 562773 493256 562779 493290
rect 562733 493218 562779 493256
rect 562733 493184 562739 493218
rect 562773 493184 562779 493218
rect 562733 493146 562779 493184
rect 562733 493112 562739 493146
rect 562773 493112 562779 493146
rect 562733 493074 562779 493112
rect 562733 493040 562739 493074
rect 562773 493040 562779 493074
rect 562733 493002 562779 493040
rect 562733 492968 562739 493002
rect 562773 492968 562779 493002
rect 562733 492930 562779 492968
rect 562733 492896 562739 492930
rect 562773 492896 562779 492930
rect 562733 492858 562779 492896
rect 562733 492824 562739 492858
rect 562773 492824 562779 492858
rect 562733 492786 562779 492824
rect 562733 492752 562739 492786
rect 562773 492752 562779 492786
rect 562733 492714 562779 492752
rect 562733 492680 562739 492714
rect 562773 492680 562779 492714
rect 562733 492642 562779 492680
rect 562733 492608 562739 492642
rect 562773 492608 562779 492642
rect 562733 492570 562779 492608
rect 562733 492536 562739 492570
rect 562773 492536 562779 492570
rect 562733 492498 562779 492536
rect 562733 492464 562739 492498
rect 562773 492464 562779 492498
rect 562733 492449 562779 492464
rect 562991 493434 563037 493449
rect 562991 493400 562997 493434
rect 563031 493400 563037 493434
rect 562991 493362 563037 493400
rect 562991 493328 562997 493362
rect 563031 493328 563037 493362
rect 562991 493290 563037 493328
rect 562991 493256 562997 493290
rect 563031 493256 563037 493290
rect 562991 493218 563037 493256
rect 562991 493184 562997 493218
rect 563031 493184 563037 493218
rect 562991 493146 563037 493184
rect 562991 493112 562997 493146
rect 563031 493112 563037 493146
rect 562991 493074 563037 493112
rect 562991 493040 562997 493074
rect 563031 493040 563037 493074
rect 562991 493002 563037 493040
rect 562991 492968 562997 493002
rect 563031 492968 563037 493002
rect 562991 492930 563037 492968
rect 562991 492896 562997 492930
rect 563031 492896 563037 492930
rect 562991 492858 563037 492896
rect 562991 492824 562997 492858
rect 563031 492824 563037 492858
rect 562991 492786 563037 492824
rect 562991 492752 562997 492786
rect 563031 492752 563037 492786
rect 562991 492714 563037 492752
rect 562991 492680 562997 492714
rect 563031 492680 563037 492714
rect 562991 492642 563037 492680
rect 562991 492608 562997 492642
rect 563031 492608 563037 492642
rect 562991 492570 563037 492608
rect 562991 492536 562997 492570
rect 563031 492536 563037 492570
rect 562991 492498 563037 492536
rect 562991 492464 562997 492498
rect 563031 492464 563037 492498
rect 562991 492449 563037 492464
rect 563249 493434 563295 493449
rect 563249 493400 563255 493434
rect 563289 493400 563295 493434
rect 563249 493362 563295 493400
rect 563249 493328 563255 493362
rect 563289 493328 563295 493362
rect 563249 493290 563295 493328
rect 563249 493256 563255 493290
rect 563289 493256 563295 493290
rect 563249 493218 563295 493256
rect 563249 493184 563255 493218
rect 563289 493184 563295 493218
rect 563249 493146 563295 493184
rect 563249 493112 563255 493146
rect 563289 493112 563295 493146
rect 563249 493074 563295 493112
rect 563249 493040 563255 493074
rect 563289 493040 563295 493074
rect 563249 493002 563295 493040
rect 563249 492968 563255 493002
rect 563289 492968 563295 493002
rect 563249 492930 563295 492968
rect 563249 492896 563255 492930
rect 563289 492896 563295 492930
rect 563249 492858 563295 492896
rect 563249 492824 563255 492858
rect 563289 492824 563295 492858
rect 563249 492786 563295 492824
rect 563249 492752 563255 492786
rect 563289 492752 563295 492786
rect 563249 492714 563295 492752
rect 563249 492680 563255 492714
rect 563289 492680 563295 492714
rect 563249 492642 563295 492680
rect 563249 492608 563255 492642
rect 563289 492608 563295 492642
rect 563249 492570 563295 492608
rect 563249 492536 563255 492570
rect 563289 492536 563295 492570
rect 563249 492498 563295 492536
rect 563249 492464 563255 492498
rect 563289 492464 563295 492498
rect 563249 492449 563295 492464
rect 563507 493434 563553 493449
rect 563507 493400 563513 493434
rect 563547 493400 563553 493434
rect 563507 493362 563553 493400
rect 563507 493328 563513 493362
rect 563547 493328 563553 493362
rect 563507 493290 563553 493328
rect 563507 493256 563513 493290
rect 563547 493256 563553 493290
rect 563507 493218 563553 493256
rect 563507 493184 563513 493218
rect 563547 493184 563553 493218
rect 563507 493146 563553 493184
rect 563507 493112 563513 493146
rect 563547 493112 563553 493146
rect 563507 493074 563553 493112
rect 563507 493040 563513 493074
rect 563547 493040 563553 493074
rect 563507 493002 563553 493040
rect 563507 492968 563513 493002
rect 563547 492968 563553 493002
rect 563507 492930 563553 492968
rect 563507 492896 563513 492930
rect 563547 492896 563553 492930
rect 563507 492858 563553 492896
rect 563507 492824 563513 492858
rect 563547 492824 563553 492858
rect 563507 492786 563553 492824
rect 563507 492752 563513 492786
rect 563547 492752 563553 492786
rect 563507 492714 563553 492752
rect 563507 492680 563513 492714
rect 563547 492680 563553 492714
rect 563507 492642 563553 492680
rect 563507 492608 563513 492642
rect 563547 492608 563553 492642
rect 563507 492570 563553 492608
rect 563507 492536 563513 492570
rect 563547 492536 563553 492570
rect 563507 492498 563553 492536
rect 563507 492464 563513 492498
rect 563547 492464 563553 492498
rect 563507 492449 563553 492464
rect 563765 493434 563811 493449
rect 563765 493400 563771 493434
rect 563805 493400 563811 493434
rect 563765 493362 563811 493400
rect 563765 493328 563771 493362
rect 563805 493328 563811 493362
rect 563765 493290 563811 493328
rect 563765 493256 563771 493290
rect 563805 493256 563811 493290
rect 563765 493218 563811 493256
rect 563765 493184 563771 493218
rect 563805 493184 563811 493218
rect 563765 493146 563811 493184
rect 563765 493112 563771 493146
rect 563805 493112 563811 493146
rect 563765 493074 563811 493112
rect 563765 493040 563771 493074
rect 563805 493040 563811 493074
rect 563765 493002 563811 493040
rect 563765 492968 563771 493002
rect 563805 492968 563811 493002
rect 563765 492930 563811 492968
rect 563765 492896 563771 492930
rect 563805 492896 563811 492930
rect 563765 492858 563811 492896
rect 563765 492824 563771 492858
rect 563805 492824 563811 492858
rect 563765 492786 563811 492824
rect 563765 492752 563771 492786
rect 563805 492752 563811 492786
rect 563765 492714 563811 492752
rect 563765 492680 563771 492714
rect 563805 492680 563811 492714
rect 563765 492642 563811 492680
rect 563765 492608 563771 492642
rect 563805 492608 563811 492642
rect 563765 492570 563811 492608
rect 563765 492536 563771 492570
rect 563805 492536 563811 492570
rect 563765 492498 563811 492536
rect 563765 492464 563771 492498
rect 563805 492464 563811 492498
rect 563765 492449 563811 492464
rect 564023 493434 564069 493449
rect 564023 493400 564029 493434
rect 564063 493400 564069 493434
rect 564023 493362 564069 493400
rect 564023 493328 564029 493362
rect 564063 493328 564069 493362
rect 564023 493290 564069 493328
rect 564023 493256 564029 493290
rect 564063 493256 564069 493290
rect 564023 493218 564069 493256
rect 564023 493184 564029 493218
rect 564063 493184 564069 493218
rect 564023 493146 564069 493184
rect 564023 493112 564029 493146
rect 564063 493112 564069 493146
rect 564023 493074 564069 493112
rect 564023 493040 564029 493074
rect 564063 493040 564069 493074
rect 564023 493002 564069 493040
rect 564023 492968 564029 493002
rect 564063 492968 564069 493002
rect 564023 492930 564069 492968
rect 564023 492896 564029 492930
rect 564063 492896 564069 492930
rect 564023 492858 564069 492896
rect 564023 492824 564029 492858
rect 564063 492824 564069 492858
rect 564023 492786 564069 492824
rect 564023 492752 564029 492786
rect 564063 492752 564069 492786
rect 564023 492714 564069 492752
rect 564023 492680 564029 492714
rect 564063 492680 564069 492714
rect 564023 492642 564069 492680
rect 564023 492608 564029 492642
rect 564063 492608 564069 492642
rect 564023 492570 564069 492608
rect 564023 492536 564029 492570
rect 564063 492536 564069 492570
rect 564023 492498 564069 492536
rect 564023 492464 564029 492498
rect 564063 492464 564069 492498
rect 564023 492449 564069 492464
rect 564281 493434 564327 493449
rect 564281 493400 564287 493434
rect 564321 493400 564327 493434
rect 564281 493362 564327 493400
rect 564281 493328 564287 493362
rect 564321 493328 564327 493362
rect 564281 493290 564327 493328
rect 564281 493256 564287 493290
rect 564321 493256 564327 493290
rect 564281 493218 564327 493256
rect 564281 493184 564287 493218
rect 564321 493184 564327 493218
rect 564281 493146 564327 493184
rect 564281 493112 564287 493146
rect 564321 493112 564327 493146
rect 564281 493074 564327 493112
rect 564281 493040 564287 493074
rect 564321 493040 564327 493074
rect 564281 493002 564327 493040
rect 564281 492968 564287 493002
rect 564321 492968 564327 493002
rect 564281 492930 564327 492968
rect 564281 492896 564287 492930
rect 564321 492896 564327 492930
rect 564281 492858 564327 492896
rect 564281 492824 564287 492858
rect 564321 492824 564327 492858
rect 564281 492786 564327 492824
rect 564281 492752 564287 492786
rect 564321 492752 564327 492786
rect 564281 492714 564327 492752
rect 564281 492680 564287 492714
rect 564321 492680 564327 492714
rect 564281 492642 564327 492680
rect 564281 492608 564287 492642
rect 564321 492608 564327 492642
rect 564281 492570 564327 492608
rect 564281 492536 564287 492570
rect 564321 492536 564327 492570
rect 564281 492498 564327 492536
rect 564281 492464 564287 492498
rect 564321 492464 564327 492498
rect 564281 492449 564327 492464
rect 564539 493434 564585 493449
rect 564539 493400 564545 493434
rect 564579 493400 564585 493434
rect 564539 493362 564585 493400
rect 564539 493328 564545 493362
rect 564579 493328 564585 493362
rect 564539 493290 564585 493328
rect 564539 493256 564545 493290
rect 564579 493256 564585 493290
rect 564539 493218 564585 493256
rect 564539 493184 564545 493218
rect 564579 493184 564585 493218
rect 564539 493146 564585 493184
rect 564539 493112 564545 493146
rect 564579 493112 564585 493146
rect 564539 493074 564585 493112
rect 564539 493040 564545 493074
rect 564579 493040 564585 493074
rect 564539 493002 564585 493040
rect 564539 492968 564545 493002
rect 564579 492968 564585 493002
rect 564539 492930 564585 492968
rect 564539 492896 564545 492930
rect 564579 492896 564585 492930
rect 564539 492858 564585 492896
rect 564539 492824 564545 492858
rect 564579 492824 564585 492858
rect 564539 492786 564585 492824
rect 564539 492752 564545 492786
rect 564579 492752 564585 492786
rect 564539 492714 564585 492752
rect 564539 492680 564545 492714
rect 564579 492680 564585 492714
rect 564539 492642 564585 492680
rect 564539 492608 564545 492642
rect 564579 492608 564585 492642
rect 564539 492570 564585 492608
rect 564539 492536 564545 492570
rect 564579 492536 564585 492570
rect 564539 492498 564585 492536
rect 564539 492464 564545 492498
rect 564579 492464 564585 492498
rect 564539 492449 564585 492464
rect 564797 493434 564843 493449
rect 564797 493400 564803 493434
rect 564837 493400 564843 493434
rect 564797 493362 564843 493400
rect 564797 493328 564803 493362
rect 564837 493328 564843 493362
rect 564797 493290 564843 493328
rect 564797 493256 564803 493290
rect 564837 493256 564843 493290
rect 564797 493218 564843 493256
rect 564797 493184 564803 493218
rect 564837 493184 564843 493218
rect 564797 493146 564843 493184
rect 564797 493112 564803 493146
rect 564837 493112 564843 493146
rect 564797 493074 564843 493112
rect 564797 493040 564803 493074
rect 564837 493040 564843 493074
rect 564797 493002 564843 493040
rect 564797 492968 564803 493002
rect 564837 492968 564843 493002
rect 564797 492930 564843 492968
rect 564797 492896 564803 492930
rect 564837 492896 564843 492930
rect 564797 492858 564843 492896
rect 564797 492824 564803 492858
rect 564837 492824 564843 492858
rect 564797 492786 564843 492824
rect 564797 492752 564803 492786
rect 564837 492752 564843 492786
rect 564797 492714 564843 492752
rect 564797 492680 564803 492714
rect 564837 492680 564843 492714
rect 564797 492642 564843 492680
rect 564797 492608 564803 492642
rect 564837 492608 564843 492642
rect 564797 492570 564843 492608
rect 564797 492536 564803 492570
rect 564837 492536 564843 492570
rect 564797 492498 564843 492536
rect 564797 492464 564803 492498
rect 564837 492464 564843 492498
rect 564797 492449 564843 492464
rect 565055 493434 565101 493449
rect 565055 493400 565061 493434
rect 565095 493400 565101 493434
rect 565055 493362 565101 493400
rect 565055 493328 565061 493362
rect 565095 493328 565101 493362
rect 565055 493290 565101 493328
rect 565055 493256 565061 493290
rect 565095 493256 565101 493290
rect 565055 493218 565101 493256
rect 565055 493184 565061 493218
rect 565095 493184 565101 493218
rect 565055 493146 565101 493184
rect 565055 493112 565061 493146
rect 565095 493112 565101 493146
rect 565055 493074 565101 493112
rect 565055 493040 565061 493074
rect 565095 493040 565101 493074
rect 565055 493002 565101 493040
rect 565055 492968 565061 493002
rect 565095 492968 565101 493002
rect 565055 492930 565101 492968
rect 565055 492896 565061 492930
rect 565095 492896 565101 492930
rect 565055 492858 565101 492896
rect 565055 492824 565061 492858
rect 565095 492824 565101 492858
rect 565055 492786 565101 492824
rect 565055 492752 565061 492786
rect 565095 492752 565101 492786
rect 565055 492714 565101 492752
rect 565055 492680 565061 492714
rect 565095 492680 565101 492714
rect 565055 492642 565101 492680
rect 565055 492608 565061 492642
rect 565095 492608 565101 492642
rect 565055 492570 565101 492608
rect 565055 492536 565061 492570
rect 565095 492536 565101 492570
rect 565055 492498 565101 492536
rect 565055 492464 565061 492498
rect 565095 492464 565101 492498
rect 565055 492449 565101 492464
rect 565313 493434 565359 493449
rect 565313 493400 565319 493434
rect 565353 493400 565359 493434
rect 565313 493362 565359 493400
rect 565313 493328 565319 493362
rect 565353 493328 565359 493362
rect 565313 493290 565359 493328
rect 565313 493256 565319 493290
rect 565353 493256 565359 493290
rect 565313 493218 565359 493256
rect 565313 493184 565319 493218
rect 565353 493184 565359 493218
rect 565313 493146 565359 493184
rect 565313 493112 565319 493146
rect 565353 493112 565359 493146
rect 565313 493074 565359 493112
rect 565313 493040 565319 493074
rect 565353 493040 565359 493074
rect 565313 493002 565359 493040
rect 565313 492968 565319 493002
rect 565353 492968 565359 493002
rect 565313 492930 565359 492968
rect 565313 492896 565319 492930
rect 565353 492896 565359 492930
rect 565313 492858 565359 492896
rect 565313 492824 565319 492858
rect 565353 492824 565359 492858
rect 565313 492786 565359 492824
rect 565313 492752 565319 492786
rect 565353 492752 565359 492786
rect 565313 492714 565359 492752
rect 565313 492680 565319 492714
rect 565353 492680 565359 492714
rect 565313 492642 565359 492680
rect 565313 492608 565319 492642
rect 565353 492608 565359 492642
rect 565313 492570 565359 492608
rect 565313 492536 565319 492570
rect 565353 492536 565359 492570
rect 565313 492498 565359 492536
rect 565313 492464 565319 492498
rect 565353 492464 565359 492498
rect 565313 492449 565359 492464
rect 565571 493434 565617 493449
rect 565571 493400 565577 493434
rect 565611 493400 565617 493434
rect 565571 493362 565617 493400
rect 565571 493328 565577 493362
rect 565611 493328 565617 493362
rect 565571 493290 565617 493328
rect 565571 493256 565577 493290
rect 565611 493256 565617 493290
rect 565571 493218 565617 493256
rect 565571 493184 565577 493218
rect 565611 493184 565617 493218
rect 565571 493146 565617 493184
rect 565571 493112 565577 493146
rect 565611 493112 565617 493146
rect 565571 493074 565617 493112
rect 565571 493040 565577 493074
rect 565611 493040 565617 493074
rect 565571 493002 565617 493040
rect 565571 492968 565577 493002
rect 565611 492968 565617 493002
rect 565571 492930 565617 492968
rect 565571 492896 565577 492930
rect 565611 492896 565617 492930
rect 565571 492858 565617 492896
rect 565571 492824 565577 492858
rect 565611 492824 565617 492858
rect 565571 492786 565617 492824
rect 565571 492752 565577 492786
rect 565611 492752 565617 492786
rect 565571 492714 565617 492752
rect 565571 492680 565577 492714
rect 565611 492680 565617 492714
rect 565571 492642 565617 492680
rect 565571 492608 565577 492642
rect 565611 492608 565617 492642
rect 565571 492570 565617 492608
rect 565571 492536 565577 492570
rect 565611 492536 565617 492570
rect 565571 492498 565617 492536
rect 565571 492464 565577 492498
rect 565611 492464 565617 492498
rect 565571 492449 565617 492464
rect 565829 493434 565875 493449
rect 565829 493400 565835 493434
rect 565869 493400 565875 493434
rect 565829 493362 565875 493400
rect 565829 493328 565835 493362
rect 565869 493328 565875 493362
rect 565829 493290 565875 493328
rect 565829 493256 565835 493290
rect 565869 493256 565875 493290
rect 565829 493218 565875 493256
rect 565829 493184 565835 493218
rect 565869 493184 565875 493218
rect 565829 493146 565875 493184
rect 565829 493112 565835 493146
rect 565869 493112 565875 493146
rect 565829 493074 565875 493112
rect 565829 493040 565835 493074
rect 565869 493040 565875 493074
rect 565829 493002 565875 493040
rect 565829 492968 565835 493002
rect 565869 492968 565875 493002
rect 565829 492930 565875 492968
rect 565829 492896 565835 492930
rect 565869 492896 565875 492930
rect 565829 492858 565875 492896
rect 565829 492824 565835 492858
rect 565869 492824 565875 492858
rect 565829 492786 565875 492824
rect 565829 492752 565835 492786
rect 565869 492752 565875 492786
rect 565829 492714 565875 492752
rect 565829 492680 565835 492714
rect 565869 492680 565875 492714
rect 565829 492642 565875 492680
rect 565829 492608 565835 492642
rect 565869 492608 565875 492642
rect 565829 492570 565875 492608
rect 565829 492536 565835 492570
rect 565869 492536 565875 492570
rect 565829 492498 565875 492536
rect 566210 492521 566418 494135
rect 573598 493667 573810 494771
rect 580860 494341 581064 494357
rect 580860 494161 580872 494341
rect 581052 494161 581064 494341
rect 580860 494145 581064 494161
rect 573598 493663 573994 493667
rect 565829 492464 565835 492498
rect 565869 492464 565875 492498
rect 565829 492449 565875 492464
rect 566048 492461 566418 492521
rect 573590 493620 580570 493663
rect 573590 493586 575255 493620
rect 575289 493586 575455 493620
rect 575489 493586 575655 493620
rect 575689 493586 575855 493620
rect 575889 493586 576055 493620
rect 576089 493586 576255 493620
rect 576289 493586 576455 493620
rect 576489 493586 576655 493620
rect 576689 493586 576855 493620
rect 576889 493586 577055 493620
rect 577089 493586 577255 493620
rect 577289 493586 577455 493620
rect 577489 493586 577655 493620
rect 577689 493586 577855 493620
rect 577889 493586 578055 493620
rect 578089 493586 578255 493620
rect 578289 493586 578455 493620
rect 578489 493586 578655 493620
rect 578689 493586 578855 493620
rect 578889 493586 579055 493620
rect 579089 493586 579255 493620
rect 579289 493586 579455 493620
rect 579489 493586 579655 493620
rect 579689 493586 579855 493620
rect 579889 493586 580055 493620
rect 580089 493586 580255 493620
rect 580289 493586 580570 493620
rect 573590 493543 580570 493586
rect 560011 492349 560500 492363
rect 559802 492313 560500 492349
rect 566048 492436 566540 492461
rect 566048 492330 566115 492436
rect 566221 492330 566540 492436
rect 566048 492313 566540 492330
rect 559802 492009 560010 492313
rect 573590 492205 573810 493543
rect 575225 493208 575271 493223
rect 575225 493174 575231 493208
rect 575265 493174 575271 493208
rect 575225 493136 575271 493174
rect 575225 493102 575231 493136
rect 575265 493102 575271 493136
rect 575225 493064 575271 493102
rect 575225 493030 575231 493064
rect 575265 493030 575271 493064
rect 575225 492992 575271 493030
rect 575225 492958 575231 492992
rect 575265 492958 575271 492992
rect 575225 492920 575271 492958
rect 575225 492886 575231 492920
rect 575265 492886 575271 492920
rect 575225 492848 575271 492886
rect 575225 492814 575231 492848
rect 575265 492814 575271 492848
rect 575225 492776 575271 492814
rect 575225 492742 575231 492776
rect 575265 492742 575271 492776
rect 575225 492704 575271 492742
rect 575225 492670 575231 492704
rect 575265 492670 575271 492704
rect 575225 492632 575271 492670
rect 575225 492598 575231 492632
rect 575265 492598 575271 492632
rect 575225 492560 575271 492598
rect 575225 492526 575231 492560
rect 575265 492526 575271 492560
rect 575225 492488 575271 492526
rect 575225 492454 575231 492488
rect 575265 492454 575271 492488
rect 575225 492416 575271 492454
rect 575225 492382 575231 492416
rect 575265 492382 575271 492416
rect 575225 492344 575271 492382
rect 575225 492310 575231 492344
rect 575265 492310 575271 492344
rect 575225 492272 575271 492310
rect 575225 492238 575231 492272
rect 575265 492238 575271 492272
rect 575225 492223 575271 492238
rect 575483 493208 575529 493223
rect 575483 493174 575489 493208
rect 575523 493174 575529 493208
rect 575483 493136 575529 493174
rect 575483 493102 575489 493136
rect 575523 493102 575529 493136
rect 575483 493064 575529 493102
rect 575483 493030 575489 493064
rect 575523 493030 575529 493064
rect 575483 492992 575529 493030
rect 575483 492958 575489 492992
rect 575523 492958 575529 492992
rect 575483 492920 575529 492958
rect 575483 492886 575489 492920
rect 575523 492886 575529 492920
rect 575483 492848 575529 492886
rect 575483 492814 575489 492848
rect 575523 492814 575529 492848
rect 575483 492776 575529 492814
rect 575483 492742 575489 492776
rect 575523 492742 575529 492776
rect 575483 492704 575529 492742
rect 575483 492670 575489 492704
rect 575523 492670 575529 492704
rect 575483 492632 575529 492670
rect 575483 492598 575489 492632
rect 575523 492598 575529 492632
rect 575483 492560 575529 492598
rect 575483 492526 575489 492560
rect 575523 492526 575529 492560
rect 575483 492488 575529 492526
rect 575483 492454 575489 492488
rect 575523 492454 575529 492488
rect 575483 492416 575529 492454
rect 575483 492382 575489 492416
rect 575523 492382 575529 492416
rect 575483 492344 575529 492382
rect 575483 492310 575489 492344
rect 575523 492310 575529 492344
rect 575483 492272 575529 492310
rect 575483 492238 575489 492272
rect 575523 492238 575529 492272
rect 575483 492223 575529 492238
rect 575741 493208 575787 493223
rect 575741 493174 575747 493208
rect 575781 493174 575787 493208
rect 575741 493136 575787 493174
rect 575741 493102 575747 493136
rect 575781 493102 575787 493136
rect 575741 493064 575787 493102
rect 575741 493030 575747 493064
rect 575781 493030 575787 493064
rect 575741 492992 575787 493030
rect 575741 492958 575747 492992
rect 575781 492958 575787 492992
rect 575741 492920 575787 492958
rect 575741 492886 575747 492920
rect 575781 492886 575787 492920
rect 575741 492848 575787 492886
rect 575741 492814 575747 492848
rect 575781 492814 575787 492848
rect 575741 492776 575787 492814
rect 575741 492742 575747 492776
rect 575781 492742 575787 492776
rect 575741 492704 575787 492742
rect 575741 492670 575747 492704
rect 575781 492670 575787 492704
rect 575741 492632 575787 492670
rect 575741 492598 575747 492632
rect 575781 492598 575787 492632
rect 575741 492560 575787 492598
rect 575741 492526 575747 492560
rect 575781 492526 575787 492560
rect 575741 492488 575787 492526
rect 575741 492454 575747 492488
rect 575781 492454 575787 492488
rect 575741 492416 575787 492454
rect 575741 492382 575747 492416
rect 575781 492382 575787 492416
rect 575741 492344 575787 492382
rect 575741 492310 575747 492344
rect 575781 492310 575787 492344
rect 575741 492272 575787 492310
rect 575741 492238 575747 492272
rect 575781 492238 575787 492272
rect 575741 492223 575787 492238
rect 575999 493208 576045 493223
rect 575999 493174 576005 493208
rect 576039 493174 576045 493208
rect 575999 493136 576045 493174
rect 575999 493102 576005 493136
rect 576039 493102 576045 493136
rect 575999 493064 576045 493102
rect 575999 493030 576005 493064
rect 576039 493030 576045 493064
rect 575999 492992 576045 493030
rect 575999 492958 576005 492992
rect 576039 492958 576045 492992
rect 575999 492920 576045 492958
rect 575999 492886 576005 492920
rect 576039 492886 576045 492920
rect 575999 492848 576045 492886
rect 575999 492814 576005 492848
rect 576039 492814 576045 492848
rect 575999 492776 576045 492814
rect 575999 492742 576005 492776
rect 576039 492742 576045 492776
rect 575999 492704 576045 492742
rect 575999 492670 576005 492704
rect 576039 492670 576045 492704
rect 575999 492632 576045 492670
rect 575999 492598 576005 492632
rect 576039 492598 576045 492632
rect 575999 492560 576045 492598
rect 575999 492526 576005 492560
rect 576039 492526 576045 492560
rect 575999 492488 576045 492526
rect 575999 492454 576005 492488
rect 576039 492454 576045 492488
rect 575999 492416 576045 492454
rect 575999 492382 576005 492416
rect 576039 492382 576045 492416
rect 575999 492344 576045 492382
rect 575999 492310 576005 492344
rect 576039 492310 576045 492344
rect 575999 492272 576045 492310
rect 575999 492238 576005 492272
rect 576039 492238 576045 492272
rect 575999 492223 576045 492238
rect 576257 493208 576303 493223
rect 576257 493174 576263 493208
rect 576297 493174 576303 493208
rect 576257 493136 576303 493174
rect 576257 493102 576263 493136
rect 576297 493102 576303 493136
rect 576257 493064 576303 493102
rect 576257 493030 576263 493064
rect 576297 493030 576303 493064
rect 576257 492992 576303 493030
rect 576257 492958 576263 492992
rect 576297 492958 576303 492992
rect 576257 492920 576303 492958
rect 576257 492886 576263 492920
rect 576297 492886 576303 492920
rect 576257 492848 576303 492886
rect 576257 492814 576263 492848
rect 576297 492814 576303 492848
rect 576257 492776 576303 492814
rect 576257 492742 576263 492776
rect 576297 492742 576303 492776
rect 576257 492704 576303 492742
rect 576257 492670 576263 492704
rect 576297 492670 576303 492704
rect 576257 492632 576303 492670
rect 576257 492598 576263 492632
rect 576297 492598 576303 492632
rect 576257 492560 576303 492598
rect 576257 492526 576263 492560
rect 576297 492526 576303 492560
rect 576257 492488 576303 492526
rect 576257 492454 576263 492488
rect 576297 492454 576303 492488
rect 576257 492416 576303 492454
rect 576257 492382 576263 492416
rect 576297 492382 576303 492416
rect 576257 492344 576303 492382
rect 576257 492310 576263 492344
rect 576297 492310 576303 492344
rect 576257 492272 576303 492310
rect 576257 492238 576263 492272
rect 576297 492238 576303 492272
rect 576257 492223 576303 492238
rect 576515 493208 576561 493223
rect 576515 493174 576521 493208
rect 576555 493174 576561 493208
rect 576515 493136 576561 493174
rect 576515 493102 576521 493136
rect 576555 493102 576561 493136
rect 576515 493064 576561 493102
rect 576515 493030 576521 493064
rect 576555 493030 576561 493064
rect 576515 492992 576561 493030
rect 576515 492958 576521 492992
rect 576555 492958 576561 492992
rect 576515 492920 576561 492958
rect 576515 492886 576521 492920
rect 576555 492886 576561 492920
rect 576515 492848 576561 492886
rect 576515 492814 576521 492848
rect 576555 492814 576561 492848
rect 576515 492776 576561 492814
rect 576515 492742 576521 492776
rect 576555 492742 576561 492776
rect 576515 492704 576561 492742
rect 576515 492670 576521 492704
rect 576555 492670 576561 492704
rect 576515 492632 576561 492670
rect 576515 492598 576521 492632
rect 576555 492598 576561 492632
rect 576515 492560 576561 492598
rect 576515 492526 576521 492560
rect 576555 492526 576561 492560
rect 576515 492488 576561 492526
rect 576515 492454 576521 492488
rect 576555 492454 576561 492488
rect 576515 492416 576561 492454
rect 576515 492382 576521 492416
rect 576555 492382 576561 492416
rect 576515 492344 576561 492382
rect 576515 492310 576521 492344
rect 576555 492310 576561 492344
rect 576515 492272 576561 492310
rect 576515 492238 576521 492272
rect 576555 492238 576561 492272
rect 576515 492223 576561 492238
rect 576773 493208 576819 493223
rect 576773 493174 576779 493208
rect 576813 493174 576819 493208
rect 576773 493136 576819 493174
rect 576773 493102 576779 493136
rect 576813 493102 576819 493136
rect 576773 493064 576819 493102
rect 576773 493030 576779 493064
rect 576813 493030 576819 493064
rect 576773 492992 576819 493030
rect 576773 492958 576779 492992
rect 576813 492958 576819 492992
rect 576773 492920 576819 492958
rect 576773 492886 576779 492920
rect 576813 492886 576819 492920
rect 576773 492848 576819 492886
rect 576773 492814 576779 492848
rect 576813 492814 576819 492848
rect 576773 492776 576819 492814
rect 576773 492742 576779 492776
rect 576813 492742 576819 492776
rect 576773 492704 576819 492742
rect 576773 492670 576779 492704
rect 576813 492670 576819 492704
rect 576773 492632 576819 492670
rect 576773 492598 576779 492632
rect 576813 492598 576819 492632
rect 576773 492560 576819 492598
rect 576773 492526 576779 492560
rect 576813 492526 576819 492560
rect 576773 492488 576819 492526
rect 576773 492454 576779 492488
rect 576813 492454 576819 492488
rect 576773 492416 576819 492454
rect 576773 492382 576779 492416
rect 576813 492382 576819 492416
rect 576773 492344 576819 492382
rect 576773 492310 576779 492344
rect 576813 492310 576819 492344
rect 576773 492272 576819 492310
rect 576773 492238 576779 492272
rect 576813 492238 576819 492272
rect 576773 492223 576819 492238
rect 577031 493208 577077 493223
rect 577031 493174 577037 493208
rect 577071 493174 577077 493208
rect 577031 493136 577077 493174
rect 577031 493102 577037 493136
rect 577071 493102 577077 493136
rect 577031 493064 577077 493102
rect 577031 493030 577037 493064
rect 577071 493030 577077 493064
rect 577031 492992 577077 493030
rect 577031 492958 577037 492992
rect 577071 492958 577077 492992
rect 577031 492920 577077 492958
rect 577031 492886 577037 492920
rect 577071 492886 577077 492920
rect 577031 492848 577077 492886
rect 577031 492814 577037 492848
rect 577071 492814 577077 492848
rect 577031 492776 577077 492814
rect 577031 492742 577037 492776
rect 577071 492742 577077 492776
rect 577031 492704 577077 492742
rect 577031 492670 577037 492704
rect 577071 492670 577077 492704
rect 577031 492632 577077 492670
rect 577031 492598 577037 492632
rect 577071 492598 577077 492632
rect 577031 492560 577077 492598
rect 577031 492526 577037 492560
rect 577071 492526 577077 492560
rect 577031 492488 577077 492526
rect 577031 492454 577037 492488
rect 577071 492454 577077 492488
rect 577031 492416 577077 492454
rect 577031 492382 577037 492416
rect 577071 492382 577077 492416
rect 577031 492344 577077 492382
rect 577031 492310 577037 492344
rect 577071 492310 577077 492344
rect 577031 492272 577077 492310
rect 577031 492238 577037 492272
rect 577071 492238 577077 492272
rect 577031 492223 577077 492238
rect 577289 493208 577335 493223
rect 577289 493174 577295 493208
rect 577329 493174 577335 493208
rect 577289 493136 577335 493174
rect 577289 493102 577295 493136
rect 577329 493102 577335 493136
rect 577289 493064 577335 493102
rect 577289 493030 577295 493064
rect 577329 493030 577335 493064
rect 577289 492992 577335 493030
rect 577289 492958 577295 492992
rect 577329 492958 577335 492992
rect 577289 492920 577335 492958
rect 577289 492886 577295 492920
rect 577329 492886 577335 492920
rect 577289 492848 577335 492886
rect 577289 492814 577295 492848
rect 577329 492814 577335 492848
rect 577289 492776 577335 492814
rect 577289 492742 577295 492776
rect 577329 492742 577335 492776
rect 577289 492704 577335 492742
rect 577289 492670 577295 492704
rect 577329 492670 577335 492704
rect 577289 492632 577335 492670
rect 577289 492598 577295 492632
rect 577329 492598 577335 492632
rect 577289 492560 577335 492598
rect 577289 492526 577295 492560
rect 577329 492526 577335 492560
rect 577289 492488 577335 492526
rect 577289 492454 577295 492488
rect 577329 492454 577335 492488
rect 577289 492416 577335 492454
rect 577289 492382 577295 492416
rect 577329 492382 577335 492416
rect 577289 492344 577335 492382
rect 577289 492310 577295 492344
rect 577329 492310 577335 492344
rect 577289 492272 577335 492310
rect 577289 492238 577295 492272
rect 577329 492238 577335 492272
rect 577289 492223 577335 492238
rect 577547 493208 577593 493223
rect 577547 493174 577553 493208
rect 577587 493174 577593 493208
rect 577547 493136 577593 493174
rect 577547 493102 577553 493136
rect 577587 493102 577593 493136
rect 577547 493064 577593 493102
rect 577547 493030 577553 493064
rect 577587 493030 577593 493064
rect 577547 492992 577593 493030
rect 577547 492958 577553 492992
rect 577587 492958 577593 492992
rect 577547 492920 577593 492958
rect 577547 492886 577553 492920
rect 577587 492886 577593 492920
rect 577547 492848 577593 492886
rect 577547 492814 577553 492848
rect 577587 492814 577593 492848
rect 577547 492776 577593 492814
rect 577547 492742 577553 492776
rect 577587 492742 577593 492776
rect 577547 492704 577593 492742
rect 577547 492670 577553 492704
rect 577587 492670 577593 492704
rect 577547 492632 577593 492670
rect 577547 492598 577553 492632
rect 577587 492598 577593 492632
rect 577547 492560 577593 492598
rect 577547 492526 577553 492560
rect 577587 492526 577593 492560
rect 577547 492488 577593 492526
rect 577547 492454 577553 492488
rect 577587 492454 577593 492488
rect 577547 492416 577593 492454
rect 577547 492382 577553 492416
rect 577587 492382 577593 492416
rect 577547 492344 577593 492382
rect 577547 492310 577553 492344
rect 577587 492310 577593 492344
rect 577547 492272 577593 492310
rect 577547 492238 577553 492272
rect 577587 492238 577593 492272
rect 577547 492223 577593 492238
rect 577805 493208 577851 493223
rect 577805 493174 577811 493208
rect 577845 493174 577851 493208
rect 577805 493136 577851 493174
rect 577805 493102 577811 493136
rect 577845 493102 577851 493136
rect 577805 493064 577851 493102
rect 577805 493030 577811 493064
rect 577845 493030 577851 493064
rect 577805 492992 577851 493030
rect 577805 492958 577811 492992
rect 577845 492958 577851 492992
rect 577805 492920 577851 492958
rect 577805 492886 577811 492920
rect 577845 492886 577851 492920
rect 577805 492848 577851 492886
rect 577805 492814 577811 492848
rect 577845 492814 577851 492848
rect 577805 492776 577851 492814
rect 577805 492742 577811 492776
rect 577845 492742 577851 492776
rect 577805 492704 577851 492742
rect 577805 492670 577811 492704
rect 577845 492670 577851 492704
rect 577805 492632 577851 492670
rect 577805 492598 577811 492632
rect 577845 492598 577851 492632
rect 577805 492560 577851 492598
rect 577805 492526 577811 492560
rect 577845 492526 577851 492560
rect 577805 492488 577851 492526
rect 577805 492454 577811 492488
rect 577845 492454 577851 492488
rect 577805 492416 577851 492454
rect 577805 492382 577811 492416
rect 577845 492382 577851 492416
rect 577805 492344 577851 492382
rect 577805 492310 577811 492344
rect 577845 492310 577851 492344
rect 577805 492272 577851 492310
rect 577805 492238 577811 492272
rect 577845 492238 577851 492272
rect 577805 492223 577851 492238
rect 578063 493208 578109 493223
rect 578063 493174 578069 493208
rect 578103 493174 578109 493208
rect 578063 493136 578109 493174
rect 578063 493102 578069 493136
rect 578103 493102 578109 493136
rect 578063 493064 578109 493102
rect 578063 493030 578069 493064
rect 578103 493030 578109 493064
rect 578063 492992 578109 493030
rect 578063 492958 578069 492992
rect 578103 492958 578109 492992
rect 578063 492920 578109 492958
rect 578063 492886 578069 492920
rect 578103 492886 578109 492920
rect 578063 492848 578109 492886
rect 578063 492814 578069 492848
rect 578103 492814 578109 492848
rect 578063 492776 578109 492814
rect 578063 492742 578069 492776
rect 578103 492742 578109 492776
rect 578063 492704 578109 492742
rect 578063 492670 578069 492704
rect 578103 492670 578109 492704
rect 578063 492632 578109 492670
rect 578063 492598 578069 492632
rect 578103 492598 578109 492632
rect 578063 492560 578109 492598
rect 578063 492526 578069 492560
rect 578103 492526 578109 492560
rect 578063 492488 578109 492526
rect 578063 492454 578069 492488
rect 578103 492454 578109 492488
rect 578063 492416 578109 492454
rect 578063 492382 578069 492416
rect 578103 492382 578109 492416
rect 578063 492344 578109 492382
rect 578063 492310 578069 492344
rect 578103 492310 578109 492344
rect 578063 492272 578109 492310
rect 578063 492238 578069 492272
rect 578103 492238 578109 492272
rect 578063 492223 578109 492238
rect 578321 493208 578367 493223
rect 578321 493174 578327 493208
rect 578361 493174 578367 493208
rect 578321 493136 578367 493174
rect 578321 493102 578327 493136
rect 578361 493102 578367 493136
rect 578321 493064 578367 493102
rect 578321 493030 578327 493064
rect 578361 493030 578367 493064
rect 578321 492992 578367 493030
rect 578321 492958 578327 492992
rect 578361 492958 578367 492992
rect 578321 492920 578367 492958
rect 578321 492886 578327 492920
rect 578361 492886 578367 492920
rect 578321 492848 578367 492886
rect 578321 492814 578327 492848
rect 578361 492814 578367 492848
rect 578321 492776 578367 492814
rect 578321 492742 578327 492776
rect 578361 492742 578367 492776
rect 578321 492704 578367 492742
rect 578321 492670 578327 492704
rect 578361 492670 578367 492704
rect 578321 492632 578367 492670
rect 578321 492598 578327 492632
rect 578361 492598 578367 492632
rect 578321 492560 578367 492598
rect 578321 492526 578327 492560
rect 578361 492526 578367 492560
rect 578321 492488 578367 492526
rect 578321 492454 578327 492488
rect 578361 492454 578367 492488
rect 578321 492416 578367 492454
rect 578321 492382 578327 492416
rect 578361 492382 578367 492416
rect 578321 492344 578367 492382
rect 578321 492310 578327 492344
rect 578361 492310 578367 492344
rect 578321 492272 578367 492310
rect 578321 492238 578327 492272
rect 578361 492238 578367 492272
rect 578321 492223 578367 492238
rect 578579 493208 578625 493223
rect 578579 493174 578585 493208
rect 578619 493174 578625 493208
rect 578579 493136 578625 493174
rect 578579 493102 578585 493136
rect 578619 493102 578625 493136
rect 578579 493064 578625 493102
rect 578579 493030 578585 493064
rect 578619 493030 578625 493064
rect 578579 492992 578625 493030
rect 578579 492958 578585 492992
rect 578619 492958 578625 492992
rect 578579 492920 578625 492958
rect 578579 492886 578585 492920
rect 578619 492886 578625 492920
rect 578579 492848 578625 492886
rect 578579 492814 578585 492848
rect 578619 492814 578625 492848
rect 578579 492776 578625 492814
rect 578579 492742 578585 492776
rect 578619 492742 578625 492776
rect 578579 492704 578625 492742
rect 578579 492670 578585 492704
rect 578619 492670 578625 492704
rect 578579 492632 578625 492670
rect 578579 492598 578585 492632
rect 578619 492598 578625 492632
rect 578579 492560 578625 492598
rect 578579 492526 578585 492560
rect 578619 492526 578625 492560
rect 578579 492488 578625 492526
rect 578579 492454 578585 492488
rect 578619 492454 578625 492488
rect 578579 492416 578625 492454
rect 578579 492382 578585 492416
rect 578619 492382 578625 492416
rect 578579 492344 578625 492382
rect 578579 492310 578585 492344
rect 578619 492310 578625 492344
rect 578579 492272 578625 492310
rect 578579 492238 578585 492272
rect 578619 492238 578625 492272
rect 578579 492223 578625 492238
rect 578837 493208 578883 493223
rect 578837 493174 578843 493208
rect 578877 493174 578883 493208
rect 578837 493136 578883 493174
rect 578837 493102 578843 493136
rect 578877 493102 578883 493136
rect 578837 493064 578883 493102
rect 578837 493030 578843 493064
rect 578877 493030 578883 493064
rect 578837 492992 578883 493030
rect 578837 492958 578843 492992
rect 578877 492958 578883 492992
rect 578837 492920 578883 492958
rect 578837 492886 578843 492920
rect 578877 492886 578883 492920
rect 578837 492848 578883 492886
rect 578837 492814 578843 492848
rect 578877 492814 578883 492848
rect 578837 492776 578883 492814
rect 578837 492742 578843 492776
rect 578877 492742 578883 492776
rect 578837 492704 578883 492742
rect 578837 492670 578843 492704
rect 578877 492670 578883 492704
rect 578837 492632 578883 492670
rect 578837 492598 578843 492632
rect 578877 492598 578883 492632
rect 578837 492560 578883 492598
rect 578837 492526 578843 492560
rect 578877 492526 578883 492560
rect 578837 492488 578883 492526
rect 578837 492454 578843 492488
rect 578877 492454 578883 492488
rect 578837 492416 578883 492454
rect 578837 492382 578843 492416
rect 578877 492382 578883 492416
rect 578837 492344 578883 492382
rect 578837 492310 578843 492344
rect 578877 492310 578883 492344
rect 578837 492272 578883 492310
rect 578837 492238 578843 492272
rect 578877 492238 578883 492272
rect 578837 492223 578883 492238
rect 579095 493208 579141 493223
rect 579095 493174 579101 493208
rect 579135 493174 579141 493208
rect 579095 493136 579141 493174
rect 579095 493102 579101 493136
rect 579135 493102 579141 493136
rect 579095 493064 579141 493102
rect 579095 493030 579101 493064
rect 579135 493030 579141 493064
rect 579095 492992 579141 493030
rect 579095 492958 579101 492992
rect 579135 492958 579141 492992
rect 579095 492920 579141 492958
rect 579095 492886 579101 492920
rect 579135 492886 579141 492920
rect 579095 492848 579141 492886
rect 579095 492814 579101 492848
rect 579135 492814 579141 492848
rect 579095 492776 579141 492814
rect 579095 492742 579101 492776
rect 579135 492742 579141 492776
rect 579095 492704 579141 492742
rect 579095 492670 579101 492704
rect 579135 492670 579141 492704
rect 579095 492632 579141 492670
rect 579095 492598 579101 492632
rect 579135 492598 579141 492632
rect 579095 492560 579141 492598
rect 579095 492526 579101 492560
rect 579135 492526 579141 492560
rect 579095 492488 579141 492526
rect 579095 492454 579101 492488
rect 579135 492454 579141 492488
rect 579095 492416 579141 492454
rect 579095 492382 579101 492416
rect 579135 492382 579141 492416
rect 579095 492344 579141 492382
rect 579095 492310 579101 492344
rect 579135 492310 579141 492344
rect 579095 492272 579141 492310
rect 579095 492238 579101 492272
rect 579135 492238 579141 492272
rect 579095 492223 579141 492238
rect 579353 493208 579399 493223
rect 579353 493174 579359 493208
rect 579393 493174 579399 493208
rect 579353 493136 579399 493174
rect 579353 493102 579359 493136
rect 579393 493102 579399 493136
rect 579353 493064 579399 493102
rect 579353 493030 579359 493064
rect 579393 493030 579399 493064
rect 579353 492992 579399 493030
rect 579353 492958 579359 492992
rect 579393 492958 579399 492992
rect 579353 492920 579399 492958
rect 579353 492886 579359 492920
rect 579393 492886 579399 492920
rect 579353 492848 579399 492886
rect 579353 492814 579359 492848
rect 579393 492814 579399 492848
rect 579353 492776 579399 492814
rect 579353 492742 579359 492776
rect 579393 492742 579399 492776
rect 579353 492704 579399 492742
rect 579353 492670 579359 492704
rect 579393 492670 579399 492704
rect 579353 492632 579399 492670
rect 579353 492598 579359 492632
rect 579393 492598 579399 492632
rect 579353 492560 579399 492598
rect 579353 492526 579359 492560
rect 579393 492526 579399 492560
rect 579353 492488 579399 492526
rect 579353 492454 579359 492488
rect 579393 492454 579399 492488
rect 579353 492416 579399 492454
rect 579353 492382 579359 492416
rect 579393 492382 579399 492416
rect 579353 492344 579399 492382
rect 579353 492310 579359 492344
rect 579393 492310 579399 492344
rect 579353 492272 579399 492310
rect 579353 492238 579359 492272
rect 579393 492238 579399 492272
rect 579353 492223 579399 492238
rect 579611 493208 579657 493223
rect 579611 493174 579617 493208
rect 579651 493174 579657 493208
rect 579611 493136 579657 493174
rect 579611 493102 579617 493136
rect 579651 493102 579657 493136
rect 579611 493064 579657 493102
rect 579611 493030 579617 493064
rect 579651 493030 579657 493064
rect 579611 492992 579657 493030
rect 579611 492958 579617 492992
rect 579651 492958 579657 492992
rect 579611 492920 579657 492958
rect 579611 492886 579617 492920
rect 579651 492886 579657 492920
rect 579611 492848 579657 492886
rect 579611 492814 579617 492848
rect 579651 492814 579657 492848
rect 579611 492776 579657 492814
rect 579611 492742 579617 492776
rect 579651 492742 579657 492776
rect 579611 492704 579657 492742
rect 579611 492670 579617 492704
rect 579651 492670 579657 492704
rect 579611 492632 579657 492670
rect 579611 492598 579617 492632
rect 579651 492598 579657 492632
rect 579611 492560 579657 492598
rect 579611 492526 579617 492560
rect 579651 492526 579657 492560
rect 579611 492488 579657 492526
rect 579611 492454 579617 492488
rect 579651 492454 579657 492488
rect 579611 492416 579657 492454
rect 579611 492382 579617 492416
rect 579651 492382 579657 492416
rect 579611 492344 579657 492382
rect 579611 492310 579617 492344
rect 579651 492310 579657 492344
rect 579611 492272 579657 492310
rect 579611 492238 579617 492272
rect 579651 492238 579657 492272
rect 579611 492223 579657 492238
rect 579869 493208 579915 493223
rect 579869 493174 579875 493208
rect 579909 493174 579915 493208
rect 579869 493136 579915 493174
rect 579869 493102 579875 493136
rect 579909 493102 579915 493136
rect 579869 493064 579915 493102
rect 579869 493030 579875 493064
rect 579909 493030 579915 493064
rect 579869 492992 579915 493030
rect 579869 492958 579875 492992
rect 579909 492958 579915 492992
rect 579869 492920 579915 492958
rect 579869 492886 579875 492920
rect 579909 492886 579915 492920
rect 579869 492848 579915 492886
rect 579869 492814 579875 492848
rect 579909 492814 579915 492848
rect 579869 492776 579915 492814
rect 579869 492742 579875 492776
rect 579909 492742 579915 492776
rect 579869 492704 579915 492742
rect 579869 492670 579875 492704
rect 579909 492670 579915 492704
rect 579869 492632 579915 492670
rect 579869 492598 579875 492632
rect 579909 492598 579915 492632
rect 579869 492560 579915 492598
rect 579869 492526 579875 492560
rect 579909 492526 579915 492560
rect 579869 492488 579915 492526
rect 579869 492454 579875 492488
rect 579909 492454 579915 492488
rect 579869 492416 579915 492454
rect 579869 492382 579875 492416
rect 579909 492382 579915 492416
rect 579869 492344 579915 492382
rect 579869 492310 579875 492344
rect 579909 492310 579915 492344
rect 579869 492272 579915 492310
rect 579869 492238 579875 492272
rect 579909 492238 579915 492272
rect 579869 492223 579915 492238
rect 580127 493208 580173 493223
rect 580127 493174 580133 493208
rect 580167 493174 580173 493208
rect 580127 493136 580173 493174
rect 580127 493102 580133 493136
rect 580167 493102 580173 493136
rect 580127 493064 580173 493102
rect 580127 493030 580133 493064
rect 580167 493030 580173 493064
rect 580127 492992 580173 493030
rect 580127 492958 580133 492992
rect 580167 492958 580173 492992
rect 580127 492920 580173 492958
rect 580127 492886 580133 492920
rect 580167 492886 580173 492920
rect 580127 492848 580173 492886
rect 580127 492814 580133 492848
rect 580167 492814 580173 492848
rect 580127 492776 580173 492814
rect 580127 492742 580133 492776
rect 580167 492742 580173 492776
rect 580127 492704 580173 492742
rect 580127 492670 580133 492704
rect 580167 492670 580173 492704
rect 580127 492632 580173 492670
rect 580127 492598 580133 492632
rect 580167 492598 580173 492632
rect 580127 492560 580173 492598
rect 580127 492526 580133 492560
rect 580167 492526 580173 492560
rect 580127 492488 580173 492526
rect 580127 492454 580133 492488
rect 580167 492454 580173 492488
rect 580127 492416 580173 492454
rect 580127 492382 580133 492416
rect 580167 492382 580173 492416
rect 580127 492344 580173 492382
rect 580127 492310 580133 492344
rect 580167 492310 580173 492344
rect 580127 492272 580173 492310
rect 580127 492238 580133 492272
rect 580167 492238 580173 492272
rect 580127 492223 580173 492238
rect 580385 493208 580431 493223
rect 580385 493174 580391 493208
rect 580425 493174 580431 493208
rect 580385 493136 580431 493174
rect 580385 493102 580391 493136
rect 580425 493102 580431 493136
rect 580385 493064 580431 493102
rect 580385 493030 580391 493064
rect 580425 493030 580431 493064
rect 580385 492992 580431 493030
rect 580385 492958 580391 492992
rect 580425 492958 580431 492992
rect 580385 492920 580431 492958
rect 580385 492886 580391 492920
rect 580425 492886 580431 492920
rect 580385 492848 580431 492886
rect 580385 492814 580391 492848
rect 580425 492814 580431 492848
rect 580385 492776 580431 492814
rect 580385 492742 580391 492776
rect 580425 492742 580431 492776
rect 580385 492704 580431 492742
rect 580385 492670 580391 492704
rect 580425 492670 580431 492704
rect 580385 492632 580431 492670
rect 580385 492598 580391 492632
rect 580425 492598 580431 492632
rect 580385 492560 580431 492598
rect 580385 492526 580391 492560
rect 580425 492526 580431 492560
rect 580385 492488 580431 492526
rect 580385 492454 580391 492488
rect 580425 492454 580431 492488
rect 580385 492416 580431 492454
rect 580385 492382 580391 492416
rect 580425 492382 580431 492416
rect 580385 492344 580431 492382
rect 580385 492310 580391 492344
rect 580425 492310 580431 492344
rect 580385 492272 580431 492310
rect 580385 492238 580391 492272
rect 580425 492238 580431 492272
rect 580385 492223 580431 492238
rect 573520 492155 573968 492205
rect 559802 491966 565978 492009
rect 559802 491932 560863 491966
rect 560897 491932 561063 491966
rect 561097 491932 561263 491966
rect 561297 491932 561463 491966
rect 561497 491932 561663 491966
rect 561697 491932 561863 491966
rect 561897 491932 562063 491966
rect 562097 491932 562263 491966
rect 562297 491932 562463 491966
rect 562497 491932 562663 491966
rect 562697 491932 562863 491966
rect 562897 491932 563063 491966
rect 563097 491932 563263 491966
rect 563297 491932 563463 491966
rect 563497 491932 563663 491966
rect 563697 491932 563863 491966
rect 563897 491932 564063 491966
rect 564097 491932 564263 491966
rect 564297 491932 564463 491966
rect 564497 491932 564663 491966
rect 564697 491932 564863 491966
rect 564897 491932 565063 491966
rect 565097 491932 565263 491966
rect 565297 491932 565463 491966
rect 565497 491932 565663 491966
rect 565697 491932 565978 491966
rect 559802 491893 565978 491932
rect 559848 491889 565978 491893
rect 573520 491911 573579 492155
rect 573887 492085 573968 492155
rect 580866 492139 581054 494145
rect 580544 492100 581054 492139
rect 573887 491958 575052 492085
rect 580544 492066 580584 492100
rect 580618 492066 581054 492100
rect 580544 492035 581054 492066
rect 580544 492033 580658 492035
rect 573887 491924 574977 491958
rect 575011 491957 575052 491958
rect 575011 491924 575048 491957
rect 573887 491911 575048 491924
rect 565740 491613 565860 491889
rect 573520 491877 575048 491911
rect 575184 491740 580570 491783
rect 575184 491706 575255 491740
rect 575289 491706 575455 491740
rect 575489 491706 575655 491740
rect 575689 491706 575855 491740
rect 575889 491706 576055 491740
rect 576089 491706 576255 491740
rect 576289 491706 576455 491740
rect 576489 491706 576655 491740
rect 576689 491706 576855 491740
rect 576889 491706 577055 491740
rect 577089 491706 577255 491740
rect 577289 491706 577455 491740
rect 577489 491706 577655 491740
rect 577689 491706 577855 491740
rect 577889 491706 578055 491740
rect 578089 491706 578255 491740
rect 578289 491706 578455 491740
rect 578489 491706 578655 491740
rect 578689 491706 578855 491740
rect 578889 491706 579055 491740
rect 579089 491706 579255 491740
rect 579289 491706 579455 491740
rect 579489 491706 579655 491740
rect 579689 491706 579855 491740
rect 579889 491706 580055 491740
rect 580089 491706 580255 491740
rect 580289 491706 580570 491740
rect 575184 491663 580570 491706
rect 575302 491613 575422 491663
rect 565740 491493 575422 491613
rect 560606 406081 573728 406201
rect 560606 404747 560726 406081
rect 566268 405485 566476 405497
rect 566260 405466 566486 405485
rect 566260 405286 566283 405466
rect 566463 405286 566486 405466
rect 566260 405267 566486 405286
rect 560600 404704 565958 404747
rect 560600 404670 560799 404704
rect 560833 404670 560999 404704
rect 561033 404670 561199 404704
rect 561233 404670 561399 404704
rect 561433 404670 561599 404704
rect 561633 404670 561799 404704
rect 561833 404670 561999 404704
rect 562033 404670 562199 404704
rect 562233 404670 562399 404704
rect 562433 404670 562599 404704
rect 562633 404670 562799 404704
rect 562833 404670 562999 404704
rect 563033 404670 563199 404704
rect 563233 404670 563399 404704
rect 563433 404670 563599 404704
rect 563633 404670 563799 404704
rect 563833 404670 563999 404704
rect 564033 404670 564199 404704
rect 564233 404670 564399 404704
rect 564433 404670 564599 404704
rect 564633 404670 564799 404704
rect 564833 404670 564999 404704
rect 565033 404670 565199 404704
rect 565233 404670 565399 404704
rect 565433 404670 565599 404704
rect 565633 404670 565958 404704
rect 560600 404627 565958 404670
rect 560605 404292 560651 404307
rect 560605 404258 560611 404292
rect 560645 404258 560651 404292
rect 560605 404220 560651 404258
rect 560605 404186 560611 404220
rect 560645 404186 560651 404220
rect 560605 404148 560651 404186
rect 560605 404114 560611 404148
rect 560645 404114 560651 404148
rect 560605 404076 560651 404114
rect 560605 404042 560611 404076
rect 560645 404042 560651 404076
rect 560605 404004 560651 404042
rect 560605 403970 560611 404004
rect 560645 403970 560651 404004
rect 560605 403932 560651 403970
rect 560605 403898 560611 403932
rect 560645 403898 560651 403932
rect 560605 403860 560651 403898
rect 560605 403826 560611 403860
rect 560645 403826 560651 403860
rect 560605 403788 560651 403826
rect 560605 403754 560611 403788
rect 560645 403754 560651 403788
rect 560605 403716 560651 403754
rect 560605 403682 560611 403716
rect 560645 403682 560651 403716
rect 560605 403644 560651 403682
rect 560605 403610 560611 403644
rect 560645 403610 560651 403644
rect 560605 403572 560651 403610
rect 560605 403538 560611 403572
rect 560645 403538 560651 403572
rect 559720 403379 560134 403501
rect 560605 403500 560651 403538
rect 560605 403466 560611 403500
rect 560645 403466 560651 403500
rect 560605 403428 560651 403466
rect 560605 403394 560611 403428
rect 560645 403394 560651 403428
rect 559720 403347 560436 403379
rect 559720 403289 559755 403347
rect 559718 403231 559755 403289
rect 559935 403327 560436 403347
rect 559935 403231 560303 403327
rect 559718 403221 560303 403231
rect 560409 403221 560436 403327
rect 560605 403356 560651 403394
rect 560605 403322 560611 403356
rect 560645 403322 560651 403356
rect 560605 403307 560651 403322
rect 560863 404292 560909 404307
rect 560863 404258 560869 404292
rect 560903 404258 560909 404292
rect 560863 404220 560909 404258
rect 560863 404186 560869 404220
rect 560903 404186 560909 404220
rect 560863 404148 560909 404186
rect 560863 404114 560869 404148
rect 560903 404114 560909 404148
rect 560863 404076 560909 404114
rect 560863 404042 560869 404076
rect 560903 404042 560909 404076
rect 560863 404004 560909 404042
rect 560863 403970 560869 404004
rect 560903 403970 560909 404004
rect 560863 403932 560909 403970
rect 560863 403898 560869 403932
rect 560903 403898 560909 403932
rect 560863 403860 560909 403898
rect 560863 403826 560869 403860
rect 560903 403826 560909 403860
rect 560863 403788 560909 403826
rect 560863 403754 560869 403788
rect 560903 403754 560909 403788
rect 560863 403716 560909 403754
rect 560863 403682 560869 403716
rect 560903 403682 560909 403716
rect 560863 403644 560909 403682
rect 560863 403610 560869 403644
rect 560903 403610 560909 403644
rect 560863 403572 560909 403610
rect 560863 403538 560869 403572
rect 560903 403538 560909 403572
rect 560863 403500 560909 403538
rect 560863 403466 560869 403500
rect 560903 403466 560909 403500
rect 560863 403428 560909 403466
rect 560863 403394 560869 403428
rect 560903 403394 560909 403428
rect 560863 403356 560909 403394
rect 560863 403322 560869 403356
rect 560903 403322 560909 403356
rect 560863 403307 560909 403322
rect 561121 404292 561167 404307
rect 561121 404258 561127 404292
rect 561161 404258 561167 404292
rect 561121 404220 561167 404258
rect 561121 404186 561127 404220
rect 561161 404186 561167 404220
rect 561121 404148 561167 404186
rect 561121 404114 561127 404148
rect 561161 404114 561167 404148
rect 561121 404076 561167 404114
rect 561121 404042 561127 404076
rect 561161 404042 561167 404076
rect 561121 404004 561167 404042
rect 561121 403970 561127 404004
rect 561161 403970 561167 404004
rect 561121 403932 561167 403970
rect 561121 403898 561127 403932
rect 561161 403898 561167 403932
rect 561121 403860 561167 403898
rect 561121 403826 561127 403860
rect 561161 403826 561167 403860
rect 561121 403788 561167 403826
rect 561121 403754 561127 403788
rect 561161 403754 561167 403788
rect 561121 403716 561167 403754
rect 561121 403682 561127 403716
rect 561161 403682 561167 403716
rect 561121 403644 561167 403682
rect 561121 403610 561127 403644
rect 561161 403610 561167 403644
rect 561121 403572 561167 403610
rect 561121 403538 561127 403572
rect 561161 403538 561167 403572
rect 561121 403500 561167 403538
rect 561121 403466 561127 403500
rect 561161 403466 561167 403500
rect 561121 403428 561167 403466
rect 561121 403394 561127 403428
rect 561161 403394 561167 403428
rect 561121 403356 561167 403394
rect 561121 403322 561127 403356
rect 561161 403322 561167 403356
rect 561121 403307 561167 403322
rect 561379 404292 561425 404307
rect 561379 404258 561385 404292
rect 561419 404258 561425 404292
rect 561379 404220 561425 404258
rect 561379 404186 561385 404220
rect 561419 404186 561425 404220
rect 561379 404148 561425 404186
rect 561379 404114 561385 404148
rect 561419 404114 561425 404148
rect 561379 404076 561425 404114
rect 561379 404042 561385 404076
rect 561419 404042 561425 404076
rect 561379 404004 561425 404042
rect 561379 403970 561385 404004
rect 561419 403970 561425 404004
rect 561379 403932 561425 403970
rect 561379 403898 561385 403932
rect 561419 403898 561425 403932
rect 561379 403860 561425 403898
rect 561379 403826 561385 403860
rect 561419 403826 561425 403860
rect 561379 403788 561425 403826
rect 561379 403754 561385 403788
rect 561419 403754 561425 403788
rect 561379 403716 561425 403754
rect 561379 403682 561385 403716
rect 561419 403682 561425 403716
rect 561379 403644 561425 403682
rect 561379 403610 561385 403644
rect 561419 403610 561425 403644
rect 561379 403572 561425 403610
rect 561379 403538 561385 403572
rect 561419 403538 561425 403572
rect 561379 403500 561425 403538
rect 561379 403466 561385 403500
rect 561419 403466 561425 403500
rect 561379 403428 561425 403466
rect 561379 403394 561385 403428
rect 561419 403394 561425 403428
rect 561379 403356 561425 403394
rect 561379 403322 561385 403356
rect 561419 403322 561425 403356
rect 561379 403307 561425 403322
rect 561637 404292 561683 404307
rect 561637 404258 561643 404292
rect 561677 404258 561683 404292
rect 561637 404220 561683 404258
rect 561637 404186 561643 404220
rect 561677 404186 561683 404220
rect 561637 404148 561683 404186
rect 561637 404114 561643 404148
rect 561677 404114 561683 404148
rect 561637 404076 561683 404114
rect 561637 404042 561643 404076
rect 561677 404042 561683 404076
rect 561637 404004 561683 404042
rect 561637 403970 561643 404004
rect 561677 403970 561683 404004
rect 561637 403932 561683 403970
rect 561637 403898 561643 403932
rect 561677 403898 561683 403932
rect 561637 403860 561683 403898
rect 561637 403826 561643 403860
rect 561677 403826 561683 403860
rect 561637 403788 561683 403826
rect 561637 403754 561643 403788
rect 561677 403754 561683 403788
rect 561637 403716 561683 403754
rect 561637 403682 561643 403716
rect 561677 403682 561683 403716
rect 561637 403644 561683 403682
rect 561637 403610 561643 403644
rect 561677 403610 561683 403644
rect 561637 403572 561683 403610
rect 561637 403538 561643 403572
rect 561677 403538 561683 403572
rect 561637 403500 561683 403538
rect 561637 403466 561643 403500
rect 561677 403466 561683 403500
rect 561637 403428 561683 403466
rect 561637 403394 561643 403428
rect 561677 403394 561683 403428
rect 561637 403356 561683 403394
rect 561637 403322 561643 403356
rect 561677 403322 561683 403356
rect 561637 403307 561683 403322
rect 561895 404292 561941 404307
rect 561895 404258 561901 404292
rect 561935 404258 561941 404292
rect 561895 404220 561941 404258
rect 561895 404186 561901 404220
rect 561935 404186 561941 404220
rect 561895 404148 561941 404186
rect 561895 404114 561901 404148
rect 561935 404114 561941 404148
rect 561895 404076 561941 404114
rect 561895 404042 561901 404076
rect 561935 404042 561941 404076
rect 561895 404004 561941 404042
rect 561895 403970 561901 404004
rect 561935 403970 561941 404004
rect 561895 403932 561941 403970
rect 561895 403898 561901 403932
rect 561935 403898 561941 403932
rect 561895 403860 561941 403898
rect 561895 403826 561901 403860
rect 561935 403826 561941 403860
rect 561895 403788 561941 403826
rect 561895 403754 561901 403788
rect 561935 403754 561941 403788
rect 561895 403716 561941 403754
rect 561895 403682 561901 403716
rect 561935 403682 561941 403716
rect 561895 403644 561941 403682
rect 561895 403610 561901 403644
rect 561935 403610 561941 403644
rect 561895 403572 561941 403610
rect 561895 403538 561901 403572
rect 561935 403538 561941 403572
rect 561895 403500 561941 403538
rect 561895 403466 561901 403500
rect 561935 403466 561941 403500
rect 561895 403428 561941 403466
rect 561895 403394 561901 403428
rect 561935 403394 561941 403428
rect 561895 403356 561941 403394
rect 561895 403322 561901 403356
rect 561935 403322 561941 403356
rect 561895 403307 561941 403322
rect 562153 404292 562199 404307
rect 562153 404258 562159 404292
rect 562193 404258 562199 404292
rect 562153 404220 562199 404258
rect 562153 404186 562159 404220
rect 562193 404186 562199 404220
rect 562153 404148 562199 404186
rect 562153 404114 562159 404148
rect 562193 404114 562199 404148
rect 562153 404076 562199 404114
rect 562153 404042 562159 404076
rect 562193 404042 562199 404076
rect 562153 404004 562199 404042
rect 562153 403970 562159 404004
rect 562193 403970 562199 404004
rect 562153 403932 562199 403970
rect 562153 403898 562159 403932
rect 562193 403898 562199 403932
rect 562153 403860 562199 403898
rect 562153 403826 562159 403860
rect 562193 403826 562199 403860
rect 562153 403788 562199 403826
rect 562153 403754 562159 403788
rect 562193 403754 562199 403788
rect 562153 403716 562199 403754
rect 562153 403682 562159 403716
rect 562193 403682 562199 403716
rect 562153 403644 562199 403682
rect 562153 403610 562159 403644
rect 562193 403610 562199 403644
rect 562153 403572 562199 403610
rect 562153 403538 562159 403572
rect 562193 403538 562199 403572
rect 562153 403500 562199 403538
rect 562153 403466 562159 403500
rect 562193 403466 562199 403500
rect 562153 403428 562199 403466
rect 562153 403394 562159 403428
rect 562193 403394 562199 403428
rect 562153 403356 562199 403394
rect 562153 403322 562159 403356
rect 562193 403322 562199 403356
rect 562153 403307 562199 403322
rect 562411 404292 562457 404307
rect 562411 404258 562417 404292
rect 562451 404258 562457 404292
rect 562411 404220 562457 404258
rect 562411 404186 562417 404220
rect 562451 404186 562457 404220
rect 562411 404148 562457 404186
rect 562411 404114 562417 404148
rect 562451 404114 562457 404148
rect 562411 404076 562457 404114
rect 562411 404042 562417 404076
rect 562451 404042 562457 404076
rect 562411 404004 562457 404042
rect 562411 403970 562417 404004
rect 562451 403970 562457 404004
rect 562411 403932 562457 403970
rect 562411 403898 562417 403932
rect 562451 403898 562457 403932
rect 562411 403860 562457 403898
rect 562411 403826 562417 403860
rect 562451 403826 562457 403860
rect 562411 403788 562457 403826
rect 562411 403754 562417 403788
rect 562451 403754 562457 403788
rect 562411 403716 562457 403754
rect 562411 403682 562417 403716
rect 562451 403682 562457 403716
rect 562411 403644 562457 403682
rect 562411 403610 562417 403644
rect 562451 403610 562457 403644
rect 562411 403572 562457 403610
rect 562411 403538 562417 403572
rect 562451 403538 562457 403572
rect 562411 403500 562457 403538
rect 562411 403466 562417 403500
rect 562451 403466 562457 403500
rect 562411 403428 562457 403466
rect 562411 403394 562417 403428
rect 562451 403394 562457 403428
rect 562411 403356 562457 403394
rect 562411 403322 562417 403356
rect 562451 403322 562457 403356
rect 562411 403307 562457 403322
rect 562669 404292 562715 404307
rect 562669 404258 562675 404292
rect 562709 404258 562715 404292
rect 562669 404220 562715 404258
rect 562669 404186 562675 404220
rect 562709 404186 562715 404220
rect 562669 404148 562715 404186
rect 562669 404114 562675 404148
rect 562709 404114 562715 404148
rect 562669 404076 562715 404114
rect 562669 404042 562675 404076
rect 562709 404042 562715 404076
rect 562669 404004 562715 404042
rect 562669 403970 562675 404004
rect 562709 403970 562715 404004
rect 562669 403932 562715 403970
rect 562669 403898 562675 403932
rect 562709 403898 562715 403932
rect 562669 403860 562715 403898
rect 562669 403826 562675 403860
rect 562709 403826 562715 403860
rect 562669 403788 562715 403826
rect 562669 403754 562675 403788
rect 562709 403754 562715 403788
rect 562669 403716 562715 403754
rect 562669 403682 562675 403716
rect 562709 403682 562715 403716
rect 562669 403644 562715 403682
rect 562669 403610 562675 403644
rect 562709 403610 562715 403644
rect 562669 403572 562715 403610
rect 562669 403538 562675 403572
rect 562709 403538 562715 403572
rect 562669 403500 562715 403538
rect 562669 403466 562675 403500
rect 562709 403466 562715 403500
rect 562669 403428 562715 403466
rect 562669 403394 562675 403428
rect 562709 403394 562715 403428
rect 562669 403356 562715 403394
rect 562669 403322 562675 403356
rect 562709 403322 562715 403356
rect 562669 403307 562715 403322
rect 562927 404292 562973 404307
rect 562927 404258 562933 404292
rect 562967 404258 562973 404292
rect 562927 404220 562973 404258
rect 562927 404186 562933 404220
rect 562967 404186 562973 404220
rect 562927 404148 562973 404186
rect 562927 404114 562933 404148
rect 562967 404114 562973 404148
rect 562927 404076 562973 404114
rect 562927 404042 562933 404076
rect 562967 404042 562973 404076
rect 562927 404004 562973 404042
rect 562927 403970 562933 404004
rect 562967 403970 562973 404004
rect 562927 403932 562973 403970
rect 562927 403898 562933 403932
rect 562967 403898 562973 403932
rect 562927 403860 562973 403898
rect 562927 403826 562933 403860
rect 562967 403826 562973 403860
rect 562927 403788 562973 403826
rect 562927 403754 562933 403788
rect 562967 403754 562973 403788
rect 562927 403716 562973 403754
rect 562927 403682 562933 403716
rect 562967 403682 562973 403716
rect 562927 403644 562973 403682
rect 562927 403610 562933 403644
rect 562967 403610 562973 403644
rect 562927 403572 562973 403610
rect 562927 403538 562933 403572
rect 562967 403538 562973 403572
rect 562927 403500 562973 403538
rect 562927 403466 562933 403500
rect 562967 403466 562973 403500
rect 562927 403428 562973 403466
rect 562927 403394 562933 403428
rect 562967 403394 562973 403428
rect 562927 403356 562973 403394
rect 562927 403322 562933 403356
rect 562967 403322 562973 403356
rect 562927 403307 562973 403322
rect 563185 404292 563231 404307
rect 563185 404258 563191 404292
rect 563225 404258 563231 404292
rect 563185 404220 563231 404258
rect 563185 404186 563191 404220
rect 563225 404186 563231 404220
rect 563185 404148 563231 404186
rect 563185 404114 563191 404148
rect 563225 404114 563231 404148
rect 563185 404076 563231 404114
rect 563185 404042 563191 404076
rect 563225 404042 563231 404076
rect 563185 404004 563231 404042
rect 563185 403970 563191 404004
rect 563225 403970 563231 404004
rect 563185 403932 563231 403970
rect 563185 403898 563191 403932
rect 563225 403898 563231 403932
rect 563185 403860 563231 403898
rect 563185 403826 563191 403860
rect 563225 403826 563231 403860
rect 563185 403788 563231 403826
rect 563185 403754 563191 403788
rect 563225 403754 563231 403788
rect 563185 403716 563231 403754
rect 563185 403682 563191 403716
rect 563225 403682 563231 403716
rect 563185 403644 563231 403682
rect 563185 403610 563191 403644
rect 563225 403610 563231 403644
rect 563185 403572 563231 403610
rect 563185 403538 563191 403572
rect 563225 403538 563231 403572
rect 563185 403500 563231 403538
rect 563185 403466 563191 403500
rect 563225 403466 563231 403500
rect 563185 403428 563231 403466
rect 563185 403394 563191 403428
rect 563225 403394 563231 403428
rect 563185 403356 563231 403394
rect 563185 403322 563191 403356
rect 563225 403322 563231 403356
rect 563185 403307 563231 403322
rect 563443 404292 563489 404307
rect 563443 404258 563449 404292
rect 563483 404258 563489 404292
rect 563443 404220 563489 404258
rect 563443 404186 563449 404220
rect 563483 404186 563489 404220
rect 563443 404148 563489 404186
rect 563443 404114 563449 404148
rect 563483 404114 563489 404148
rect 563443 404076 563489 404114
rect 563443 404042 563449 404076
rect 563483 404042 563489 404076
rect 563443 404004 563489 404042
rect 563443 403970 563449 404004
rect 563483 403970 563489 404004
rect 563443 403932 563489 403970
rect 563443 403898 563449 403932
rect 563483 403898 563489 403932
rect 563443 403860 563489 403898
rect 563443 403826 563449 403860
rect 563483 403826 563489 403860
rect 563443 403788 563489 403826
rect 563443 403754 563449 403788
rect 563483 403754 563489 403788
rect 563443 403716 563489 403754
rect 563443 403682 563449 403716
rect 563483 403682 563489 403716
rect 563443 403644 563489 403682
rect 563443 403610 563449 403644
rect 563483 403610 563489 403644
rect 563443 403572 563489 403610
rect 563443 403538 563449 403572
rect 563483 403538 563489 403572
rect 563443 403500 563489 403538
rect 563443 403466 563449 403500
rect 563483 403466 563489 403500
rect 563443 403428 563489 403466
rect 563443 403394 563449 403428
rect 563483 403394 563489 403428
rect 563443 403356 563489 403394
rect 563443 403322 563449 403356
rect 563483 403322 563489 403356
rect 563443 403307 563489 403322
rect 563701 404292 563747 404307
rect 563701 404258 563707 404292
rect 563741 404258 563747 404292
rect 563701 404220 563747 404258
rect 563701 404186 563707 404220
rect 563741 404186 563747 404220
rect 563701 404148 563747 404186
rect 563701 404114 563707 404148
rect 563741 404114 563747 404148
rect 563701 404076 563747 404114
rect 563701 404042 563707 404076
rect 563741 404042 563747 404076
rect 563701 404004 563747 404042
rect 563701 403970 563707 404004
rect 563741 403970 563747 404004
rect 563701 403932 563747 403970
rect 563701 403898 563707 403932
rect 563741 403898 563747 403932
rect 563701 403860 563747 403898
rect 563701 403826 563707 403860
rect 563741 403826 563747 403860
rect 563701 403788 563747 403826
rect 563701 403754 563707 403788
rect 563741 403754 563747 403788
rect 563701 403716 563747 403754
rect 563701 403682 563707 403716
rect 563741 403682 563747 403716
rect 563701 403644 563747 403682
rect 563701 403610 563707 403644
rect 563741 403610 563747 403644
rect 563701 403572 563747 403610
rect 563701 403538 563707 403572
rect 563741 403538 563747 403572
rect 563701 403500 563747 403538
rect 563701 403466 563707 403500
rect 563741 403466 563747 403500
rect 563701 403428 563747 403466
rect 563701 403394 563707 403428
rect 563741 403394 563747 403428
rect 563701 403356 563747 403394
rect 563701 403322 563707 403356
rect 563741 403322 563747 403356
rect 563701 403307 563747 403322
rect 563959 404292 564005 404307
rect 563959 404258 563965 404292
rect 563999 404258 564005 404292
rect 563959 404220 564005 404258
rect 563959 404186 563965 404220
rect 563999 404186 564005 404220
rect 563959 404148 564005 404186
rect 563959 404114 563965 404148
rect 563999 404114 564005 404148
rect 563959 404076 564005 404114
rect 563959 404042 563965 404076
rect 563999 404042 564005 404076
rect 563959 404004 564005 404042
rect 563959 403970 563965 404004
rect 563999 403970 564005 404004
rect 563959 403932 564005 403970
rect 563959 403898 563965 403932
rect 563999 403898 564005 403932
rect 563959 403860 564005 403898
rect 563959 403826 563965 403860
rect 563999 403826 564005 403860
rect 563959 403788 564005 403826
rect 563959 403754 563965 403788
rect 563999 403754 564005 403788
rect 563959 403716 564005 403754
rect 563959 403682 563965 403716
rect 563999 403682 564005 403716
rect 563959 403644 564005 403682
rect 563959 403610 563965 403644
rect 563999 403610 564005 403644
rect 563959 403572 564005 403610
rect 563959 403538 563965 403572
rect 563999 403538 564005 403572
rect 563959 403500 564005 403538
rect 563959 403466 563965 403500
rect 563999 403466 564005 403500
rect 563959 403428 564005 403466
rect 563959 403394 563965 403428
rect 563999 403394 564005 403428
rect 563959 403356 564005 403394
rect 563959 403322 563965 403356
rect 563999 403322 564005 403356
rect 563959 403307 564005 403322
rect 564217 404292 564263 404307
rect 564217 404258 564223 404292
rect 564257 404258 564263 404292
rect 564217 404220 564263 404258
rect 564217 404186 564223 404220
rect 564257 404186 564263 404220
rect 564217 404148 564263 404186
rect 564217 404114 564223 404148
rect 564257 404114 564263 404148
rect 564217 404076 564263 404114
rect 564217 404042 564223 404076
rect 564257 404042 564263 404076
rect 564217 404004 564263 404042
rect 564217 403970 564223 404004
rect 564257 403970 564263 404004
rect 564217 403932 564263 403970
rect 564217 403898 564223 403932
rect 564257 403898 564263 403932
rect 564217 403860 564263 403898
rect 564217 403826 564223 403860
rect 564257 403826 564263 403860
rect 564217 403788 564263 403826
rect 564217 403754 564223 403788
rect 564257 403754 564263 403788
rect 564217 403716 564263 403754
rect 564217 403682 564223 403716
rect 564257 403682 564263 403716
rect 564217 403644 564263 403682
rect 564217 403610 564223 403644
rect 564257 403610 564263 403644
rect 564217 403572 564263 403610
rect 564217 403538 564223 403572
rect 564257 403538 564263 403572
rect 564217 403500 564263 403538
rect 564217 403466 564223 403500
rect 564257 403466 564263 403500
rect 564217 403428 564263 403466
rect 564217 403394 564223 403428
rect 564257 403394 564263 403428
rect 564217 403356 564263 403394
rect 564217 403322 564223 403356
rect 564257 403322 564263 403356
rect 564217 403307 564263 403322
rect 564475 404292 564521 404307
rect 564475 404258 564481 404292
rect 564515 404258 564521 404292
rect 564475 404220 564521 404258
rect 564475 404186 564481 404220
rect 564515 404186 564521 404220
rect 564475 404148 564521 404186
rect 564475 404114 564481 404148
rect 564515 404114 564521 404148
rect 564475 404076 564521 404114
rect 564475 404042 564481 404076
rect 564515 404042 564521 404076
rect 564475 404004 564521 404042
rect 564475 403970 564481 404004
rect 564515 403970 564521 404004
rect 564475 403932 564521 403970
rect 564475 403898 564481 403932
rect 564515 403898 564521 403932
rect 564475 403860 564521 403898
rect 564475 403826 564481 403860
rect 564515 403826 564521 403860
rect 564475 403788 564521 403826
rect 564475 403754 564481 403788
rect 564515 403754 564521 403788
rect 564475 403716 564521 403754
rect 564475 403682 564481 403716
rect 564515 403682 564521 403716
rect 564475 403644 564521 403682
rect 564475 403610 564481 403644
rect 564515 403610 564521 403644
rect 564475 403572 564521 403610
rect 564475 403538 564481 403572
rect 564515 403538 564521 403572
rect 564475 403500 564521 403538
rect 564475 403466 564481 403500
rect 564515 403466 564521 403500
rect 564475 403428 564521 403466
rect 564475 403394 564481 403428
rect 564515 403394 564521 403428
rect 564475 403356 564521 403394
rect 564475 403322 564481 403356
rect 564515 403322 564521 403356
rect 564475 403307 564521 403322
rect 564733 404292 564779 404307
rect 564733 404258 564739 404292
rect 564773 404258 564779 404292
rect 564733 404220 564779 404258
rect 564733 404186 564739 404220
rect 564773 404186 564779 404220
rect 564733 404148 564779 404186
rect 564733 404114 564739 404148
rect 564773 404114 564779 404148
rect 564733 404076 564779 404114
rect 564733 404042 564739 404076
rect 564773 404042 564779 404076
rect 564733 404004 564779 404042
rect 564733 403970 564739 404004
rect 564773 403970 564779 404004
rect 564733 403932 564779 403970
rect 564733 403898 564739 403932
rect 564773 403898 564779 403932
rect 564733 403860 564779 403898
rect 564733 403826 564739 403860
rect 564773 403826 564779 403860
rect 564733 403788 564779 403826
rect 564733 403754 564739 403788
rect 564773 403754 564779 403788
rect 564733 403716 564779 403754
rect 564733 403682 564739 403716
rect 564773 403682 564779 403716
rect 564733 403644 564779 403682
rect 564733 403610 564739 403644
rect 564773 403610 564779 403644
rect 564733 403572 564779 403610
rect 564733 403538 564739 403572
rect 564773 403538 564779 403572
rect 564733 403500 564779 403538
rect 564733 403466 564739 403500
rect 564773 403466 564779 403500
rect 564733 403428 564779 403466
rect 564733 403394 564739 403428
rect 564773 403394 564779 403428
rect 564733 403356 564779 403394
rect 564733 403322 564739 403356
rect 564773 403322 564779 403356
rect 564733 403307 564779 403322
rect 564991 404292 565037 404307
rect 564991 404258 564997 404292
rect 565031 404258 565037 404292
rect 564991 404220 565037 404258
rect 564991 404186 564997 404220
rect 565031 404186 565037 404220
rect 564991 404148 565037 404186
rect 564991 404114 564997 404148
rect 565031 404114 565037 404148
rect 564991 404076 565037 404114
rect 564991 404042 564997 404076
rect 565031 404042 565037 404076
rect 564991 404004 565037 404042
rect 564991 403970 564997 404004
rect 565031 403970 565037 404004
rect 564991 403932 565037 403970
rect 564991 403898 564997 403932
rect 565031 403898 565037 403932
rect 564991 403860 565037 403898
rect 564991 403826 564997 403860
rect 565031 403826 565037 403860
rect 564991 403788 565037 403826
rect 564991 403754 564997 403788
rect 565031 403754 565037 403788
rect 564991 403716 565037 403754
rect 564991 403682 564997 403716
rect 565031 403682 565037 403716
rect 564991 403644 565037 403682
rect 564991 403610 564997 403644
rect 565031 403610 565037 403644
rect 564991 403572 565037 403610
rect 564991 403538 564997 403572
rect 565031 403538 565037 403572
rect 564991 403500 565037 403538
rect 564991 403466 564997 403500
rect 565031 403466 565037 403500
rect 564991 403428 565037 403466
rect 564991 403394 564997 403428
rect 565031 403394 565037 403428
rect 564991 403356 565037 403394
rect 564991 403322 564997 403356
rect 565031 403322 565037 403356
rect 564991 403307 565037 403322
rect 565249 404292 565295 404307
rect 565249 404258 565255 404292
rect 565289 404258 565295 404292
rect 565249 404220 565295 404258
rect 565249 404186 565255 404220
rect 565289 404186 565295 404220
rect 565249 404148 565295 404186
rect 565249 404114 565255 404148
rect 565289 404114 565295 404148
rect 565249 404076 565295 404114
rect 565249 404042 565255 404076
rect 565289 404042 565295 404076
rect 565249 404004 565295 404042
rect 565249 403970 565255 404004
rect 565289 403970 565295 404004
rect 565249 403932 565295 403970
rect 565249 403898 565255 403932
rect 565289 403898 565295 403932
rect 565249 403860 565295 403898
rect 565249 403826 565255 403860
rect 565289 403826 565295 403860
rect 565249 403788 565295 403826
rect 565249 403754 565255 403788
rect 565289 403754 565295 403788
rect 565249 403716 565295 403754
rect 565249 403682 565255 403716
rect 565289 403682 565295 403716
rect 565249 403644 565295 403682
rect 565249 403610 565255 403644
rect 565289 403610 565295 403644
rect 565249 403572 565295 403610
rect 565249 403538 565255 403572
rect 565289 403538 565295 403572
rect 565249 403500 565295 403538
rect 565249 403466 565255 403500
rect 565289 403466 565295 403500
rect 565249 403428 565295 403466
rect 565249 403394 565255 403428
rect 565289 403394 565295 403428
rect 565249 403356 565295 403394
rect 565249 403322 565255 403356
rect 565289 403322 565295 403356
rect 565249 403307 565295 403322
rect 565507 404292 565553 404307
rect 565507 404258 565513 404292
rect 565547 404258 565553 404292
rect 565507 404220 565553 404258
rect 565507 404186 565513 404220
rect 565547 404186 565553 404220
rect 565507 404148 565553 404186
rect 565507 404114 565513 404148
rect 565547 404114 565553 404148
rect 565507 404076 565553 404114
rect 565507 404042 565513 404076
rect 565547 404042 565553 404076
rect 565507 404004 565553 404042
rect 565507 403970 565513 404004
rect 565547 403970 565553 404004
rect 565507 403932 565553 403970
rect 565507 403898 565513 403932
rect 565547 403898 565553 403932
rect 565507 403860 565553 403898
rect 565507 403826 565513 403860
rect 565547 403826 565553 403860
rect 565507 403788 565553 403826
rect 565507 403754 565513 403788
rect 565547 403754 565553 403788
rect 565507 403716 565553 403754
rect 565507 403682 565513 403716
rect 565547 403682 565553 403716
rect 565507 403644 565553 403682
rect 565507 403610 565513 403644
rect 565547 403610 565553 403644
rect 565507 403572 565553 403610
rect 565507 403538 565513 403572
rect 565547 403538 565553 403572
rect 565507 403500 565553 403538
rect 565507 403466 565513 403500
rect 565547 403466 565553 403500
rect 565507 403428 565553 403466
rect 565507 403394 565513 403428
rect 565547 403394 565553 403428
rect 565507 403356 565553 403394
rect 565507 403322 565513 403356
rect 565547 403322 565553 403356
rect 565507 403307 565553 403322
rect 565765 404292 565811 404307
rect 565765 404258 565771 404292
rect 565805 404258 565811 404292
rect 565765 404220 565811 404258
rect 565765 404186 565771 404220
rect 565805 404186 565811 404220
rect 565765 404148 565811 404186
rect 565765 404114 565771 404148
rect 565805 404114 565811 404148
rect 565765 404076 565811 404114
rect 565765 404042 565771 404076
rect 565805 404042 565811 404076
rect 565765 404004 565811 404042
rect 565765 403970 565771 404004
rect 565805 403970 565811 404004
rect 565765 403932 565811 403970
rect 565765 403898 565771 403932
rect 565805 403898 565811 403932
rect 565765 403860 565811 403898
rect 565765 403826 565771 403860
rect 565805 403826 565811 403860
rect 565765 403788 565811 403826
rect 565765 403754 565771 403788
rect 565805 403754 565811 403788
rect 565765 403716 565811 403754
rect 565765 403682 565771 403716
rect 565805 403682 565811 403716
rect 565765 403644 565811 403682
rect 565765 403610 565771 403644
rect 565805 403610 565811 403644
rect 565765 403572 565811 403610
rect 565765 403538 565771 403572
rect 565805 403538 565811 403572
rect 565765 403500 565811 403538
rect 565765 403466 565771 403500
rect 565805 403466 565811 403500
rect 565765 403428 565811 403466
rect 565765 403394 565771 403428
rect 565805 403394 565811 403428
rect 565765 403356 565811 403394
rect 565765 403322 565771 403356
rect 565805 403322 565811 403356
rect 565765 403307 565811 403322
rect 566268 403319 566476 405267
rect 573526 404883 573728 406081
rect 580090 405411 580194 405429
rect 580078 405382 580206 405411
rect 580078 405330 580116 405382
rect 580168 405330 580206 405382
rect 580078 405301 580206 405330
rect 573526 404681 574915 404883
rect 559718 403171 560436 403221
rect 566008 403294 566476 403319
rect 566008 403188 566051 403294
rect 566157 403188 566476 403294
rect 566008 403171 566476 403188
rect 573450 403244 573826 403262
rect 559718 402867 560160 403171
rect 573450 402962 573462 403244
rect 573824 403086 573834 403244
rect 580090 403116 580194 405301
rect 573824 402962 574370 403086
rect 573450 402958 574370 402962
rect 559718 402824 574946 402867
rect 559718 402790 560799 402824
rect 560833 402790 560999 402824
rect 561033 402790 561199 402824
rect 561233 402790 561399 402824
rect 561433 402790 561599 402824
rect 561633 402790 561799 402824
rect 561833 402790 561999 402824
rect 562033 402790 562199 402824
rect 562233 402790 562399 402824
rect 562433 402790 562599 402824
rect 562633 402790 562799 402824
rect 562833 402790 562999 402824
rect 563033 402790 563199 402824
rect 563233 402790 563399 402824
rect 563433 402790 563599 402824
rect 563633 402790 563799 402824
rect 563833 402790 563999 402824
rect 564033 402790 564199 402824
rect 564233 402790 564399 402824
rect 564433 402790 564599 402824
rect 564633 402790 564799 402824
rect 564833 402790 564999 402824
rect 565033 402790 565199 402824
rect 565233 402790 565399 402824
rect 565433 402790 565599 402824
rect 565633 402790 574946 402824
rect 559718 402747 574946 402790
rect 565750 360473 573810 360593
rect 565750 359429 565870 360473
rect 566284 359987 566508 360011
rect 566278 359981 566524 359987
rect 566278 359801 566311 359981
rect 566491 359801 566524 359981
rect 566278 359795 566524 359801
rect 560556 359386 565870 359429
rect 560556 359352 560755 359386
rect 560789 359352 560955 359386
rect 560989 359352 561155 359386
rect 561189 359352 561355 359386
rect 561389 359352 561555 359386
rect 561589 359352 561755 359386
rect 561789 359352 561955 359386
rect 561989 359352 562155 359386
rect 562189 359352 562355 359386
rect 562389 359352 562555 359386
rect 562589 359352 562755 359386
rect 562789 359352 562955 359386
rect 562989 359352 563155 359386
rect 563189 359352 563355 359386
rect 563389 359352 563555 359386
rect 563589 359352 563755 359386
rect 563789 359352 563955 359386
rect 563989 359352 564155 359386
rect 564189 359352 564355 359386
rect 564389 359352 564555 359386
rect 564589 359352 564755 359386
rect 564789 359352 564955 359386
rect 564989 359352 565155 359386
rect 565189 359352 565355 359386
rect 565389 359352 565555 359386
rect 565589 359352 565870 359386
rect 560556 359309 565870 359352
rect 560561 358974 560607 358989
rect 560561 358940 560567 358974
rect 560601 358940 560607 358974
rect 560561 358902 560607 358940
rect 560561 358868 560567 358902
rect 560601 358868 560607 358902
rect 560561 358830 560607 358868
rect 560561 358796 560567 358830
rect 560601 358796 560607 358830
rect 560561 358758 560607 358796
rect 560561 358724 560567 358758
rect 560601 358724 560607 358758
rect 560561 358686 560607 358724
rect 560561 358652 560567 358686
rect 560601 358652 560607 358686
rect 560561 358614 560607 358652
rect 560561 358580 560567 358614
rect 560601 358580 560607 358614
rect 560561 358542 560607 358580
rect 560561 358508 560567 358542
rect 560601 358508 560607 358542
rect 560561 358470 560607 358508
rect 560561 358436 560567 358470
rect 560601 358436 560607 358470
rect 560561 358398 560607 358436
rect 560561 358364 560567 358398
rect 560601 358364 560607 358398
rect 560561 358326 560607 358364
rect 560561 358292 560567 358326
rect 560601 358292 560607 358326
rect 560561 358254 560607 358292
rect 560561 358220 560567 358254
rect 560601 358220 560607 358254
rect 560561 358182 560607 358220
rect 560561 358148 560567 358182
rect 560601 358148 560607 358182
rect 560561 358110 560607 358148
rect 560561 358076 560567 358110
rect 560601 358076 560607 358110
rect 559716 358047 560392 358061
rect 559716 357867 559740 358047
rect 559920 358009 560392 358047
rect 559920 357903 560259 358009
rect 560365 357903 560392 358009
rect 560561 358038 560607 358076
rect 560561 358004 560567 358038
rect 560601 358004 560607 358038
rect 560561 357989 560607 358004
rect 560819 358974 560865 358989
rect 560819 358940 560825 358974
rect 560859 358940 560865 358974
rect 560819 358902 560865 358940
rect 560819 358868 560825 358902
rect 560859 358868 560865 358902
rect 560819 358830 560865 358868
rect 560819 358796 560825 358830
rect 560859 358796 560865 358830
rect 560819 358758 560865 358796
rect 560819 358724 560825 358758
rect 560859 358724 560865 358758
rect 560819 358686 560865 358724
rect 560819 358652 560825 358686
rect 560859 358652 560865 358686
rect 560819 358614 560865 358652
rect 560819 358580 560825 358614
rect 560859 358580 560865 358614
rect 560819 358542 560865 358580
rect 560819 358508 560825 358542
rect 560859 358508 560865 358542
rect 560819 358470 560865 358508
rect 560819 358436 560825 358470
rect 560859 358436 560865 358470
rect 560819 358398 560865 358436
rect 560819 358364 560825 358398
rect 560859 358364 560865 358398
rect 560819 358326 560865 358364
rect 560819 358292 560825 358326
rect 560859 358292 560865 358326
rect 560819 358254 560865 358292
rect 560819 358220 560825 358254
rect 560859 358220 560865 358254
rect 560819 358182 560865 358220
rect 560819 358148 560825 358182
rect 560859 358148 560865 358182
rect 560819 358110 560865 358148
rect 560819 358076 560825 358110
rect 560859 358076 560865 358110
rect 560819 358038 560865 358076
rect 560819 358004 560825 358038
rect 560859 358004 560865 358038
rect 560819 357989 560865 358004
rect 561077 358974 561123 358989
rect 561077 358940 561083 358974
rect 561117 358940 561123 358974
rect 561077 358902 561123 358940
rect 561077 358868 561083 358902
rect 561117 358868 561123 358902
rect 561077 358830 561123 358868
rect 561077 358796 561083 358830
rect 561117 358796 561123 358830
rect 561077 358758 561123 358796
rect 561077 358724 561083 358758
rect 561117 358724 561123 358758
rect 561077 358686 561123 358724
rect 561077 358652 561083 358686
rect 561117 358652 561123 358686
rect 561077 358614 561123 358652
rect 561077 358580 561083 358614
rect 561117 358580 561123 358614
rect 561077 358542 561123 358580
rect 561077 358508 561083 358542
rect 561117 358508 561123 358542
rect 561077 358470 561123 358508
rect 561077 358436 561083 358470
rect 561117 358436 561123 358470
rect 561077 358398 561123 358436
rect 561077 358364 561083 358398
rect 561117 358364 561123 358398
rect 561077 358326 561123 358364
rect 561077 358292 561083 358326
rect 561117 358292 561123 358326
rect 561077 358254 561123 358292
rect 561077 358220 561083 358254
rect 561117 358220 561123 358254
rect 561077 358182 561123 358220
rect 561077 358148 561083 358182
rect 561117 358148 561123 358182
rect 561077 358110 561123 358148
rect 561077 358076 561083 358110
rect 561117 358076 561123 358110
rect 561077 358038 561123 358076
rect 561077 358004 561083 358038
rect 561117 358004 561123 358038
rect 561077 357989 561123 358004
rect 561335 358974 561381 358989
rect 561335 358940 561341 358974
rect 561375 358940 561381 358974
rect 561335 358902 561381 358940
rect 561335 358868 561341 358902
rect 561375 358868 561381 358902
rect 561335 358830 561381 358868
rect 561335 358796 561341 358830
rect 561375 358796 561381 358830
rect 561335 358758 561381 358796
rect 561335 358724 561341 358758
rect 561375 358724 561381 358758
rect 561335 358686 561381 358724
rect 561335 358652 561341 358686
rect 561375 358652 561381 358686
rect 561335 358614 561381 358652
rect 561335 358580 561341 358614
rect 561375 358580 561381 358614
rect 561335 358542 561381 358580
rect 561335 358508 561341 358542
rect 561375 358508 561381 358542
rect 561335 358470 561381 358508
rect 561335 358436 561341 358470
rect 561375 358436 561381 358470
rect 561335 358398 561381 358436
rect 561335 358364 561341 358398
rect 561375 358364 561381 358398
rect 561335 358326 561381 358364
rect 561335 358292 561341 358326
rect 561375 358292 561381 358326
rect 561335 358254 561381 358292
rect 561335 358220 561341 358254
rect 561375 358220 561381 358254
rect 561335 358182 561381 358220
rect 561335 358148 561341 358182
rect 561375 358148 561381 358182
rect 561335 358110 561381 358148
rect 561335 358076 561341 358110
rect 561375 358076 561381 358110
rect 561335 358038 561381 358076
rect 561335 358004 561341 358038
rect 561375 358004 561381 358038
rect 561335 357989 561381 358004
rect 561593 358974 561639 358989
rect 561593 358940 561599 358974
rect 561633 358940 561639 358974
rect 561593 358902 561639 358940
rect 561593 358868 561599 358902
rect 561633 358868 561639 358902
rect 561593 358830 561639 358868
rect 561593 358796 561599 358830
rect 561633 358796 561639 358830
rect 561593 358758 561639 358796
rect 561593 358724 561599 358758
rect 561633 358724 561639 358758
rect 561593 358686 561639 358724
rect 561593 358652 561599 358686
rect 561633 358652 561639 358686
rect 561593 358614 561639 358652
rect 561593 358580 561599 358614
rect 561633 358580 561639 358614
rect 561593 358542 561639 358580
rect 561593 358508 561599 358542
rect 561633 358508 561639 358542
rect 561593 358470 561639 358508
rect 561593 358436 561599 358470
rect 561633 358436 561639 358470
rect 561593 358398 561639 358436
rect 561593 358364 561599 358398
rect 561633 358364 561639 358398
rect 561593 358326 561639 358364
rect 561593 358292 561599 358326
rect 561633 358292 561639 358326
rect 561593 358254 561639 358292
rect 561593 358220 561599 358254
rect 561633 358220 561639 358254
rect 561593 358182 561639 358220
rect 561593 358148 561599 358182
rect 561633 358148 561639 358182
rect 561593 358110 561639 358148
rect 561593 358076 561599 358110
rect 561633 358076 561639 358110
rect 561593 358038 561639 358076
rect 561593 358004 561599 358038
rect 561633 358004 561639 358038
rect 561593 357989 561639 358004
rect 561851 358974 561897 358989
rect 561851 358940 561857 358974
rect 561891 358940 561897 358974
rect 561851 358902 561897 358940
rect 561851 358868 561857 358902
rect 561891 358868 561897 358902
rect 561851 358830 561897 358868
rect 561851 358796 561857 358830
rect 561891 358796 561897 358830
rect 561851 358758 561897 358796
rect 561851 358724 561857 358758
rect 561891 358724 561897 358758
rect 561851 358686 561897 358724
rect 561851 358652 561857 358686
rect 561891 358652 561897 358686
rect 561851 358614 561897 358652
rect 561851 358580 561857 358614
rect 561891 358580 561897 358614
rect 561851 358542 561897 358580
rect 561851 358508 561857 358542
rect 561891 358508 561897 358542
rect 561851 358470 561897 358508
rect 561851 358436 561857 358470
rect 561891 358436 561897 358470
rect 561851 358398 561897 358436
rect 561851 358364 561857 358398
rect 561891 358364 561897 358398
rect 561851 358326 561897 358364
rect 561851 358292 561857 358326
rect 561891 358292 561897 358326
rect 561851 358254 561897 358292
rect 561851 358220 561857 358254
rect 561891 358220 561897 358254
rect 561851 358182 561897 358220
rect 561851 358148 561857 358182
rect 561891 358148 561897 358182
rect 561851 358110 561897 358148
rect 561851 358076 561857 358110
rect 561891 358076 561897 358110
rect 561851 358038 561897 358076
rect 561851 358004 561857 358038
rect 561891 358004 561897 358038
rect 561851 357989 561897 358004
rect 562109 358974 562155 358989
rect 562109 358940 562115 358974
rect 562149 358940 562155 358974
rect 562109 358902 562155 358940
rect 562109 358868 562115 358902
rect 562149 358868 562155 358902
rect 562109 358830 562155 358868
rect 562109 358796 562115 358830
rect 562149 358796 562155 358830
rect 562109 358758 562155 358796
rect 562109 358724 562115 358758
rect 562149 358724 562155 358758
rect 562109 358686 562155 358724
rect 562109 358652 562115 358686
rect 562149 358652 562155 358686
rect 562109 358614 562155 358652
rect 562109 358580 562115 358614
rect 562149 358580 562155 358614
rect 562109 358542 562155 358580
rect 562109 358508 562115 358542
rect 562149 358508 562155 358542
rect 562109 358470 562155 358508
rect 562109 358436 562115 358470
rect 562149 358436 562155 358470
rect 562109 358398 562155 358436
rect 562109 358364 562115 358398
rect 562149 358364 562155 358398
rect 562109 358326 562155 358364
rect 562109 358292 562115 358326
rect 562149 358292 562155 358326
rect 562109 358254 562155 358292
rect 562109 358220 562115 358254
rect 562149 358220 562155 358254
rect 562109 358182 562155 358220
rect 562109 358148 562115 358182
rect 562149 358148 562155 358182
rect 562109 358110 562155 358148
rect 562109 358076 562115 358110
rect 562149 358076 562155 358110
rect 562109 358038 562155 358076
rect 562109 358004 562115 358038
rect 562149 358004 562155 358038
rect 562109 357989 562155 358004
rect 562367 358974 562413 358989
rect 562367 358940 562373 358974
rect 562407 358940 562413 358974
rect 562367 358902 562413 358940
rect 562367 358868 562373 358902
rect 562407 358868 562413 358902
rect 562367 358830 562413 358868
rect 562367 358796 562373 358830
rect 562407 358796 562413 358830
rect 562367 358758 562413 358796
rect 562367 358724 562373 358758
rect 562407 358724 562413 358758
rect 562367 358686 562413 358724
rect 562367 358652 562373 358686
rect 562407 358652 562413 358686
rect 562367 358614 562413 358652
rect 562367 358580 562373 358614
rect 562407 358580 562413 358614
rect 562367 358542 562413 358580
rect 562367 358508 562373 358542
rect 562407 358508 562413 358542
rect 562367 358470 562413 358508
rect 562367 358436 562373 358470
rect 562407 358436 562413 358470
rect 562367 358398 562413 358436
rect 562367 358364 562373 358398
rect 562407 358364 562413 358398
rect 562367 358326 562413 358364
rect 562367 358292 562373 358326
rect 562407 358292 562413 358326
rect 562367 358254 562413 358292
rect 562367 358220 562373 358254
rect 562407 358220 562413 358254
rect 562367 358182 562413 358220
rect 562367 358148 562373 358182
rect 562407 358148 562413 358182
rect 562367 358110 562413 358148
rect 562367 358076 562373 358110
rect 562407 358076 562413 358110
rect 562367 358038 562413 358076
rect 562367 358004 562373 358038
rect 562407 358004 562413 358038
rect 562367 357989 562413 358004
rect 562625 358974 562671 358989
rect 562625 358940 562631 358974
rect 562665 358940 562671 358974
rect 562625 358902 562671 358940
rect 562625 358868 562631 358902
rect 562665 358868 562671 358902
rect 562625 358830 562671 358868
rect 562625 358796 562631 358830
rect 562665 358796 562671 358830
rect 562625 358758 562671 358796
rect 562625 358724 562631 358758
rect 562665 358724 562671 358758
rect 562625 358686 562671 358724
rect 562625 358652 562631 358686
rect 562665 358652 562671 358686
rect 562625 358614 562671 358652
rect 562625 358580 562631 358614
rect 562665 358580 562671 358614
rect 562625 358542 562671 358580
rect 562625 358508 562631 358542
rect 562665 358508 562671 358542
rect 562625 358470 562671 358508
rect 562625 358436 562631 358470
rect 562665 358436 562671 358470
rect 562625 358398 562671 358436
rect 562625 358364 562631 358398
rect 562665 358364 562671 358398
rect 562625 358326 562671 358364
rect 562625 358292 562631 358326
rect 562665 358292 562671 358326
rect 562625 358254 562671 358292
rect 562625 358220 562631 358254
rect 562665 358220 562671 358254
rect 562625 358182 562671 358220
rect 562625 358148 562631 358182
rect 562665 358148 562671 358182
rect 562625 358110 562671 358148
rect 562625 358076 562631 358110
rect 562665 358076 562671 358110
rect 562625 358038 562671 358076
rect 562625 358004 562631 358038
rect 562665 358004 562671 358038
rect 562625 357989 562671 358004
rect 562883 358974 562929 358989
rect 562883 358940 562889 358974
rect 562923 358940 562929 358974
rect 562883 358902 562929 358940
rect 562883 358868 562889 358902
rect 562923 358868 562929 358902
rect 562883 358830 562929 358868
rect 562883 358796 562889 358830
rect 562923 358796 562929 358830
rect 562883 358758 562929 358796
rect 562883 358724 562889 358758
rect 562923 358724 562929 358758
rect 562883 358686 562929 358724
rect 562883 358652 562889 358686
rect 562923 358652 562929 358686
rect 562883 358614 562929 358652
rect 562883 358580 562889 358614
rect 562923 358580 562929 358614
rect 562883 358542 562929 358580
rect 562883 358508 562889 358542
rect 562923 358508 562929 358542
rect 562883 358470 562929 358508
rect 562883 358436 562889 358470
rect 562923 358436 562929 358470
rect 562883 358398 562929 358436
rect 562883 358364 562889 358398
rect 562923 358364 562929 358398
rect 562883 358326 562929 358364
rect 562883 358292 562889 358326
rect 562923 358292 562929 358326
rect 562883 358254 562929 358292
rect 562883 358220 562889 358254
rect 562923 358220 562929 358254
rect 562883 358182 562929 358220
rect 562883 358148 562889 358182
rect 562923 358148 562929 358182
rect 562883 358110 562929 358148
rect 562883 358076 562889 358110
rect 562923 358076 562929 358110
rect 562883 358038 562929 358076
rect 562883 358004 562889 358038
rect 562923 358004 562929 358038
rect 562883 357989 562929 358004
rect 563141 358974 563187 358989
rect 563141 358940 563147 358974
rect 563181 358940 563187 358974
rect 563141 358902 563187 358940
rect 563141 358868 563147 358902
rect 563181 358868 563187 358902
rect 563141 358830 563187 358868
rect 563141 358796 563147 358830
rect 563181 358796 563187 358830
rect 563141 358758 563187 358796
rect 563141 358724 563147 358758
rect 563181 358724 563187 358758
rect 563141 358686 563187 358724
rect 563141 358652 563147 358686
rect 563181 358652 563187 358686
rect 563141 358614 563187 358652
rect 563141 358580 563147 358614
rect 563181 358580 563187 358614
rect 563141 358542 563187 358580
rect 563141 358508 563147 358542
rect 563181 358508 563187 358542
rect 563141 358470 563187 358508
rect 563141 358436 563147 358470
rect 563181 358436 563187 358470
rect 563141 358398 563187 358436
rect 563141 358364 563147 358398
rect 563181 358364 563187 358398
rect 563141 358326 563187 358364
rect 563141 358292 563147 358326
rect 563181 358292 563187 358326
rect 563141 358254 563187 358292
rect 563141 358220 563147 358254
rect 563181 358220 563187 358254
rect 563141 358182 563187 358220
rect 563141 358148 563147 358182
rect 563181 358148 563187 358182
rect 563141 358110 563187 358148
rect 563141 358076 563147 358110
rect 563181 358076 563187 358110
rect 563141 358038 563187 358076
rect 563141 358004 563147 358038
rect 563181 358004 563187 358038
rect 563141 357989 563187 358004
rect 563399 358974 563445 358989
rect 563399 358940 563405 358974
rect 563439 358940 563445 358974
rect 563399 358902 563445 358940
rect 563399 358868 563405 358902
rect 563439 358868 563445 358902
rect 563399 358830 563445 358868
rect 563399 358796 563405 358830
rect 563439 358796 563445 358830
rect 563399 358758 563445 358796
rect 563399 358724 563405 358758
rect 563439 358724 563445 358758
rect 563399 358686 563445 358724
rect 563399 358652 563405 358686
rect 563439 358652 563445 358686
rect 563399 358614 563445 358652
rect 563399 358580 563405 358614
rect 563439 358580 563445 358614
rect 563399 358542 563445 358580
rect 563399 358508 563405 358542
rect 563439 358508 563445 358542
rect 563399 358470 563445 358508
rect 563399 358436 563405 358470
rect 563439 358436 563445 358470
rect 563399 358398 563445 358436
rect 563399 358364 563405 358398
rect 563439 358364 563445 358398
rect 563399 358326 563445 358364
rect 563399 358292 563405 358326
rect 563439 358292 563445 358326
rect 563399 358254 563445 358292
rect 563399 358220 563405 358254
rect 563439 358220 563445 358254
rect 563399 358182 563445 358220
rect 563399 358148 563405 358182
rect 563439 358148 563445 358182
rect 563399 358110 563445 358148
rect 563399 358076 563405 358110
rect 563439 358076 563445 358110
rect 563399 358038 563445 358076
rect 563399 358004 563405 358038
rect 563439 358004 563445 358038
rect 563399 357989 563445 358004
rect 563657 358974 563703 358989
rect 563657 358940 563663 358974
rect 563697 358940 563703 358974
rect 563657 358902 563703 358940
rect 563657 358868 563663 358902
rect 563697 358868 563703 358902
rect 563657 358830 563703 358868
rect 563657 358796 563663 358830
rect 563697 358796 563703 358830
rect 563657 358758 563703 358796
rect 563657 358724 563663 358758
rect 563697 358724 563703 358758
rect 563657 358686 563703 358724
rect 563657 358652 563663 358686
rect 563697 358652 563703 358686
rect 563657 358614 563703 358652
rect 563657 358580 563663 358614
rect 563697 358580 563703 358614
rect 563657 358542 563703 358580
rect 563657 358508 563663 358542
rect 563697 358508 563703 358542
rect 563657 358470 563703 358508
rect 563657 358436 563663 358470
rect 563697 358436 563703 358470
rect 563657 358398 563703 358436
rect 563657 358364 563663 358398
rect 563697 358364 563703 358398
rect 563657 358326 563703 358364
rect 563657 358292 563663 358326
rect 563697 358292 563703 358326
rect 563657 358254 563703 358292
rect 563657 358220 563663 358254
rect 563697 358220 563703 358254
rect 563657 358182 563703 358220
rect 563657 358148 563663 358182
rect 563697 358148 563703 358182
rect 563657 358110 563703 358148
rect 563657 358076 563663 358110
rect 563697 358076 563703 358110
rect 563657 358038 563703 358076
rect 563657 358004 563663 358038
rect 563697 358004 563703 358038
rect 563657 357989 563703 358004
rect 563915 358974 563961 358989
rect 563915 358940 563921 358974
rect 563955 358940 563961 358974
rect 563915 358902 563961 358940
rect 563915 358868 563921 358902
rect 563955 358868 563961 358902
rect 563915 358830 563961 358868
rect 563915 358796 563921 358830
rect 563955 358796 563961 358830
rect 563915 358758 563961 358796
rect 563915 358724 563921 358758
rect 563955 358724 563961 358758
rect 563915 358686 563961 358724
rect 563915 358652 563921 358686
rect 563955 358652 563961 358686
rect 563915 358614 563961 358652
rect 563915 358580 563921 358614
rect 563955 358580 563961 358614
rect 563915 358542 563961 358580
rect 563915 358508 563921 358542
rect 563955 358508 563961 358542
rect 563915 358470 563961 358508
rect 563915 358436 563921 358470
rect 563955 358436 563961 358470
rect 563915 358398 563961 358436
rect 563915 358364 563921 358398
rect 563955 358364 563961 358398
rect 563915 358326 563961 358364
rect 563915 358292 563921 358326
rect 563955 358292 563961 358326
rect 563915 358254 563961 358292
rect 563915 358220 563921 358254
rect 563955 358220 563961 358254
rect 563915 358182 563961 358220
rect 563915 358148 563921 358182
rect 563955 358148 563961 358182
rect 563915 358110 563961 358148
rect 563915 358076 563921 358110
rect 563955 358076 563961 358110
rect 563915 358038 563961 358076
rect 563915 358004 563921 358038
rect 563955 358004 563961 358038
rect 563915 357989 563961 358004
rect 564173 358974 564219 358989
rect 564173 358940 564179 358974
rect 564213 358940 564219 358974
rect 564173 358902 564219 358940
rect 564173 358868 564179 358902
rect 564213 358868 564219 358902
rect 564173 358830 564219 358868
rect 564173 358796 564179 358830
rect 564213 358796 564219 358830
rect 564173 358758 564219 358796
rect 564173 358724 564179 358758
rect 564213 358724 564219 358758
rect 564173 358686 564219 358724
rect 564173 358652 564179 358686
rect 564213 358652 564219 358686
rect 564173 358614 564219 358652
rect 564173 358580 564179 358614
rect 564213 358580 564219 358614
rect 564173 358542 564219 358580
rect 564173 358508 564179 358542
rect 564213 358508 564219 358542
rect 564173 358470 564219 358508
rect 564173 358436 564179 358470
rect 564213 358436 564219 358470
rect 564173 358398 564219 358436
rect 564173 358364 564179 358398
rect 564213 358364 564219 358398
rect 564173 358326 564219 358364
rect 564173 358292 564179 358326
rect 564213 358292 564219 358326
rect 564173 358254 564219 358292
rect 564173 358220 564179 358254
rect 564213 358220 564219 358254
rect 564173 358182 564219 358220
rect 564173 358148 564179 358182
rect 564213 358148 564219 358182
rect 564173 358110 564219 358148
rect 564173 358076 564179 358110
rect 564213 358076 564219 358110
rect 564173 358038 564219 358076
rect 564173 358004 564179 358038
rect 564213 358004 564219 358038
rect 564173 357989 564219 358004
rect 564431 358974 564477 358989
rect 564431 358940 564437 358974
rect 564471 358940 564477 358974
rect 564431 358902 564477 358940
rect 564431 358868 564437 358902
rect 564471 358868 564477 358902
rect 564431 358830 564477 358868
rect 564431 358796 564437 358830
rect 564471 358796 564477 358830
rect 564431 358758 564477 358796
rect 564431 358724 564437 358758
rect 564471 358724 564477 358758
rect 564431 358686 564477 358724
rect 564431 358652 564437 358686
rect 564471 358652 564477 358686
rect 564431 358614 564477 358652
rect 564431 358580 564437 358614
rect 564471 358580 564477 358614
rect 564431 358542 564477 358580
rect 564431 358508 564437 358542
rect 564471 358508 564477 358542
rect 564431 358470 564477 358508
rect 564431 358436 564437 358470
rect 564471 358436 564477 358470
rect 564431 358398 564477 358436
rect 564431 358364 564437 358398
rect 564471 358364 564477 358398
rect 564431 358326 564477 358364
rect 564431 358292 564437 358326
rect 564471 358292 564477 358326
rect 564431 358254 564477 358292
rect 564431 358220 564437 358254
rect 564471 358220 564477 358254
rect 564431 358182 564477 358220
rect 564431 358148 564437 358182
rect 564471 358148 564477 358182
rect 564431 358110 564477 358148
rect 564431 358076 564437 358110
rect 564471 358076 564477 358110
rect 564431 358038 564477 358076
rect 564431 358004 564437 358038
rect 564471 358004 564477 358038
rect 564431 357989 564477 358004
rect 564689 358974 564735 358989
rect 564689 358940 564695 358974
rect 564729 358940 564735 358974
rect 564689 358902 564735 358940
rect 564689 358868 564695 358902
rect 564729 358868 564735 358902
rect 564689 358830 564735 358868
rect 564689 358796 564695 358830
rect 564729 358796 564735 358830
rect 564689 358758 564735 358796
rect 564689 358724 564695 358758
rect 564729 358724 564735 358758
rect 564689 358686 564735 358724
rect 564689 358652 564695 358686
rect 564729 358652 564735 358686
rect 564689 358614 564735 358652
rect 564689 358580 564695 358614
rect 564729 358580 564735 358614
rect 564689 358542 564735 358580
rect 564689 358508 564695 358542
rect 564729 358508 564735 358542
rect 564689 358470 564735 358508
rect 564689 358436 564695 358470
rect 564729 358436 564735 358470
rect 564689 358398 564735 358436
rect 564689 358364 564695 358398
rect 564729 358364 564735 358398
rect 564689 358326 564735 358364
rect 564689 358292 564695 358326
rect 564729 358292 564735 358326
rect 564689 358254 564735 358292
rect 564689 358220 564695 358254
rect 564729 358220 564735 358254
rect 564689 358182 564735 358220
rect 564689 358148 564695 358182
rect 564729 358148 564735 358182
rect 564689 358110 564735 358148
rect 564689 358076 564695 358110
rect 564729 358076 564735 358110
rect 564689 358038 564735 358076
rect 564689 358004 564695 358038
rect 564729 358004 564735 358038
rect 564689 357989 564735 358004
rect 564947 358974 564993 358989
rect 564947 358940 564953 358974
rect 564987 358940 564993 358974
rect 564947 358902 564993 358940
rect 564947 358868 564953 358902
rect 564987 358868 564993 358902
rect 564947 358830 564993 358868
rect 564947 358796 564953 358830
rect 564987 358796 564993 358830
rect 564947 358758 564993 358796
rect 564947 358724 564953 358758
rect 564987 358724 564993 358758
rect 564947 358686 564993 358724
rect 564947 358652 564953 358686
rect 564987 358652 564993 358686
rect 564947 358614 564993 358652
rect 564947 358580 564953 358614
rect 564987 358580 564993 358614
rect 564947 358542 564993 358580
rect 564947 358508 564953 358542
rect 564987 358508 564993 358542
rect 564947 358470 564993 358508
rect 564947 358436 564953 358470
rect 564987 358436 564993 358470
rect 564947 358398 564993 358436
rect 564947 358364 564953 358398
rect 564987 358364 564993 358398
rect 564947 358326 564993 358364
rect 564947 358292 564953 358326
rect 564987 358292 564993 358326
rect 564947 358254 564993 358292
rect 564947 358220 564953 358254
rect 564987 358220 564993 358254
rect 564947 358182 564993 358220
rect 564947 358148 564953 358182
rect 564987 358148 564993 358182
rect 564947 358110 564993 358148
rect 564947 358076 564953 358110
rect 564987 358076 564993 358110
rect 564947 358038 564993 358076
rect 564947 358004 564953 358038
rect 564987 358004 564993 358038
rect 564947 357989 564993 358004
rect 565205 358974 565251 358989
rect 565205 358940 565211 358974
rect 565245 358940 565251 358974
rect 565205 358902 565251 358940
rect 565205 358868 565211 358902
rect 565245 358868 565251 358902
rect 565205 358830 565251 358868
rect 565205 358796 565211 358830
rect 565245 358796 565251 358830
rect 565205 358758 565251 358796
rect 565205 358724 565211 358758
rect 565245 358724 565251 358758
rect 565205 358686 565251 358724
rect 565205 358652 565211 358686
rect 565245 358652 565251 358686
rect 565205 358614 565251 358652
rect 565205 358580 565211 358614
rect 565245 358580 565251 358614
rect 565205 358542 565251 358580
rect 565205 358508 565211 358542
rect 565245 358508 565251 358542
rect 565205 358470 565251 358508
rect 565205 358436 565211 358470
rect 565245 358436 565251 358470
rect 565205 358398 565251 358436
rect 565205 358364 565211 358398
rect 565245 358364 565251 358398
rect 565205 358326 565251 358364
rect 565205 358292 565211 358326
rect 565245 358292 565251 358326
rect 565205 358254 565251 358292
rect 565205 358220 565211 358254
rect 565245 358220 565251 358254
rect 565205 358182 565251 358220
rect 565205 358148 565211 358182
rect 565245 358148 565251 358182
rect 565205 358110 565251 358148
rect 565205 358076 565211 358110
rect 565245 358076 565251 358110
rect 565205 358038 565251 358076
rect 565205 358004 565211 358038
rect 565245 358004 565251 358038
rect 565205 357989 565251 358004
rect 565463 358974 565509 358989
rect 565463 358940 565469 358974
rect 565503 358940 565509 358974
rect 565463 358902 565509 358940
rect 565463 358868 565469 358902
rect 565503 358868 565509 358902
rect 565463 358830 565509 358868
rect 565463 358796 565469 358830
rect 565503 358796 565509 358830
rect 565463 358758 565509 358796
rect 565463 358724 565469 358758
rect 565503 358724 565509 358758
rect 565463 358686 565509 358724
rect 565463 358652 565469 358686
rect 565503 358652 565509 358686
rect 565463 358614 565509 358652
rect 565463 358580 565469 358614
rect 565503 358580 565509 358614
rect 565463 358542 565509 358580
rect 565463 358508 565469 358542
rect 565503 358508 565509 358542
rect 565463 358470 565509 358508
rect 565463 358436 565469 358470
rect 565503 358436 565509 358470
rect 565463 358398 565509 358436
rect 565463 358364 565469 358398
rect 565503 358364 565509 358398
rect 565463 358326 565509 358364
rect 565463 358292 565469 358326
rect 565503 358292 565509 358326
rect 565463 358254 565509 358292
rect 565463 358220 565469 358254
rect 565503 358220 565509 358254
rect 565463 358182 565509 358220
rect 565463 358148 565469 358182
rect 565503 358148 565509 358182
rect 565463 358110 565509 358148
rect 565463 358076 565469 358110
rect 565503 358076 565509 358110
rect 565463 358038 565509 358076
rect 565463 358004 565469 358038
rect 565503 358004 565509 358038
rect 565463 357989 565509 358004
rect 565721 358974 565767 358989
rect 565721 358940 565727 358974
rect 565761 358940 565767 358974
rect 565721 358902 565767 358940
rect 565721 358868 565727 358902
rect 565761 358868 565767 358902
rect 565721 358830 565767 358868
rect 565721 358796 565727 358830
rect 565761 358796 565767 358830
rect 565721 358758 565767 358796
rect 565721 358724 565727 358758
rect 565761 358724 565767 358758
rect 565721 358686 565767 358724
rect 565721 358652 565727 358686
rect 565761 358652 565767 358686
rect 565721 358614 565767 358652
rect 565721 358580 565727 358614
rect 565761 358580 565767 358614
rect 565721 358542 565767 358580
rect 565721 358508 565727 358542
rect 565761 358508 565767 358542
rect 565721 358470 565767 358508
rect 565721 358436 565727 358470
rect 565761 358436 565767 358470
rect 565721 358398 565767 358436
rect 565721 358364 565727 358398
rect 565761 358364 565767 358398
rect 565721 358326 565767 358364
rect 565721 358292 565727 358326
rect 565761 358292 565767 358326
rect 565721 358254 565767 358292
rect 565721 358220 565727 358254
rect 565761 358220 565767 358254
rect 565721 358182 565767 358220
rect 565721 358148 565727 358182
rect 565761 358148 565767 358182
rect 565721 358110 565767 358148
rect 565721 358076 565727 358110
rect 565761 358076 565767 358110
rect 565721 358038 565767 358076
rect 565721 358004 565727 358038
rect 565761 358004 565767 358038
rect 565721 357989 565767 358004
rect 566284 358001 566508 359795
rect 573602 359359 573810 360473
rect 580266 359915 580370 359943
rect 580256 359913 580382 359915
rect 580256 359861 580293 359913
rect 580345 359861 580382 359913
rect 580256 359849 580382 359861
rect 580256 359797 580293 359849
rect 580345 359797 580382 359849
rect 580256 359795 580382 359797
rect 573602 359316 580044 359359
rect 573602 359282 574729 359316
rect 574763 359282 574929 359316
rect 574963 359282 575129 359316
rect 575163 359282 575329 359316
rect 575363 359282 575529 359316
rect 575563 359282 575729 359316
rect 575763 359282 575929 359316
rect 575963 359282 576129 359316
rect 576163 359282 576329 359316
rect 576363 359282 576529 359316
rect 576563 359282 576729 359316
rect 576763 359282 576929 359316
rect 576963 359282 577129 359316
rect 577163 359282 577329 359316
rect 577363 359282 577529 359316
rect 577563 359282 577729 359316
rect 577763 359282 577929 359316
rect 577963 359282 578129 359316
rect 578163 359282 578329 359316
rect 578363 359282 578529 359316
rect 578563 359282 578729 359316
rect 578763 359282 578929 359316
rect 578963 359282 579129 359316
rect 579163 359282 579329 359316
rect 579363 359282 579529 359316
rect 579563 359282 579729 359316
rect 579763 359282 580044 359316
rect 573602 359265 580044 359282
rect 559920 357867 560392 357903
rect 559716 357853 560392 357867
rect 565964 357976 566508 358001
rect 565964 357870 566007 357976
rect 566113 357870 566508 357976
rect 573604 359239 580044 359265
rect 573604 357974 573842 359239
rect 565964 357855 566508 357870
rect 573523 357968 573842 357974
rect 574699 358904 574745 358919
rect 574699 358870 574705 358904
rect 574739 358870 574745 358904
rect 574699 358832 574745 358870
rect 574699 358798 574705 358832
rect 574739 358798 574745 358832
rect 574699 358760 574745 358798
rect 574699 358726 574705 358760
rect 574739 358726 574745 358760
rect 574699 358688 574745 358726
rect 574699 358654 574705 358688
rect 574739 358654 574745 358688
rect 574699 358616 574745 358654
rect 574699 358582 574705 358616
rect 574739 358582 574745 358616
rect 574699 358544 574745 358582
rect 574699 358510 574705 358544
rect 574739 358510 574745 358544
rect 574699 358472 574745 358510
rect 574699 358438 574705 358472
rect 574739 358438 574745 358472
rect 574699 358400 574745 358438
rect 574699 358366 574705 358400
rect 574739 358366 574745 358400
rect 574699 358328 574745 358366
rect 574699 358294 574705 358328
rect 574739 358294 574745 358328
rect 574699 358256 574745 358294
rect 574699 358222 574705 358256
rect 574739 358222 574745 358256
rect 574699 358184 574745 358222
rect 574699 358150 574705 358184
rect 574739 358150 574745 358184
rect 574699 358112 574745 358150
rect 574699 358078 574705 358112
rect 574739 358078 574745 358112
rect 574699 358040 574745 358078
rect 574699 358006 574705 358040
rect 574739 358006 574745 358040
rect 574699 357968 574745 358006
rect 573523 357920 573925 357968
rect 565964 357853 566432 357855
rect 559746 357549 559942 357853
rect 573523 357612 573569 357920
rect 573877 357819 573925 357920
rect 574699 357934 574705 357968
rect 574739 357934 574745 357968
rect 574699 357919 574745 357934
rect 574957 358904 575003 358919
rect 574957 358870 574963 358904
rect 574997 358870 575003 358904
rect 574957 358832 575003 358870
rect 574957 358798 574963 358832
rect 574997 358798 575003 358832
rect 574957 358760 575003 358798
rect 574957 358726 574963 358760
rect 574997 358726 575003 358760
rect 574957 358688 575003 358726
rect 574957 358654 574963 358688
rect 574997 358654 575003 358688
rect 574957 358616 575003 358654
rect 574957 358582 574963 358616
rect 574997 358582 575003 358616
rect 574957 358544 575003 358582
rect 574957 358510 574963 358544
rect 574997 358510 575003 358544
rect 574957 358472 575003 358510
rect 574957 358438 574963 358472
rect 574997 358438 575003 358472
rect 574957 358400 575003 358438
rect 574957 358366 574963 358400
rect 574997 358366 575003 358400
rect 574957 358328 575003 358366
rect 574957 358294 574963 358328
rect 574997 358294 575003 358328
rect 574957 358256 575003 358294
rect 574957 358222 574963 358256
rect 574997 358222 575003 358256
rect 574957 358184 575003 358222
rect 574957 358150 574963 358184
rect 574997 358150 575003 358184
rect 574957 358112 575003 358150
rect 574957 358078 574963 358112
rect 574997 358078 575003 358112
rect 574957 358040 575003 358078
rect 574957 358006 574963 358040
rect 574997 358006 575003 358040
rect 574957 357968 575003 358006
rect 574957 357934 574963 357968
rect 574997 357934 575003 357968
rect 574957 357919 575003 357934
rect 575215 358904 575261 358919
rect 575215 358870 575221 358904
rect 575255 358870 575261 358904
rect 575215 358832 575261 358870
rect 575215 358798 575221 358832
rect 575255 358798 575261 358832
rect 575215 358760 575261 358798
rect 575215 358726 575221 358760
rect 575255 358726 575261 358760
rect 575215 358688 575261 358726
rect 575215 358654 575221 358688
rect 575255 358654 575261 358688
rect 575215 358616 575261 358654
rect 575215 358582 575221 358616
rect 575255 358582 575261 358616
rect 575215 358544 575261 358582
rect 575215 358510 575221 358544
rect 575255 358510 575261 358544
rect 575215 358472 575261 358510
rect 575215 358438 575221 358472
rect 575255 358438 575261 358472
rect 575215 358400 575261 358438
rect 575215 358366 575221 358400
rect 575255 358366 575261 358400
rect 575215 358328 575261 358366
rect 575215 358294 575221 358328
rect 575255 358294 575261 358328
rect 575215 358256 575261 358294
rect 575215 358222 575221 358256
rect 575255 358222 575261 358256
rect 575215 358184 575261 358222
rect 575215 358150 575221 358184
rect 575255 358150 575261 358184
rect 575215 358112 575261 358150
rect 575215 358078 575221 358112
rect 575255 358078 575261 358112
rect 575215 358040 575261 358078
rect 575215 358006 575221 358040
rect 575255 358006 575261 358040
rect 575215 357968 575261 358006
rect 575215 357934 575221 357968
rect 575255 357934 575261 357968
rect 575215 357919 575261 357934
rect 575473 358904 575519 358919
rect 575473 358870 575479 358904
rect 575513 358870 575519 358904
rect 575473 358832 575519 358870
rect 575473 358798 575479 358832
rect 575513 358798 575519 358832
rect 575473 358760 575519 358798
rect 575473 358726 575479 358760
rect 575513 358726 575519 358760
rect 575473 358688 575519 358726
rect 575473 358654 575479 358688
rect 575513 358654 575519 358688
rect 575473 358616 575519 358654
rect 575473 358582 575479 358616
rect 575513 358582 575519 358616
rect 575473 358544 575519 358582
rect 575473 358510 575479 358544
rect 575513 358510 575519 358544
rect 575473 358472 575519 358510
rect 575473 358438 575479 358472
rect 575513 358438 575519 358472
rect 575473 358400 575519 358438
rect 575473 358366 575479 358400
rect 575513 358366 575519 358400
rect 575473 358328 575519 358366
rect 575473 358294 575479 358328
rect 575513 358294 575519 358328
rect 575473 358256 575519 358294
rect 575473 358222 575479 358256
rect 575513 358222 575519 358256
rect 575473 358184 575519 358222
rect 575473 358150 575479 358184
rect 575513 358150 575519 358184
rect 575473 358112 575519 358150
rect 575473 358078 575479 358112
rect 575513 358078 575519 358112
rect 575473 358040 575519 358078
rect 575473 358006 575479 358040
rect 575513 358006 575519 358040
rect 575473 357968 575519 358006
rect 575473 357934 575479 357968
rect 575513 357934 575519 357968
rect 575473 357919 575519 357934
rect 575731 358904 575777 358919
rect 575731 358870 575737 358904
rect 575771 358870 575777 358904
rect 575731 358832 575777 358870
rect 575731 358798 575737 358832
rect 575771 358798 575777 358832
rect 575731 358760 575777 358798
rect 575731 358726 575737 358760
rect 575771 358726 575777 358760
rect 575731 358688 575777 358726
rect 575731 358654 575737 358688
rect 575771 358654 575777 358688
rect 575731 358616 575777 358654
rect 575731 358582 575737 358616
rect 575771 358582 575777 358616
rect 575731 358544 575777 358582
rect 575731 358510 575737 358544
rect 575771 358510 575777 358544
rect 575731 358472 575777 358510
rect 575731 358438 575737 358472
rect 575771 358438 575777 358472
rect 575731 358400 575777 358438
rect 575731 358366 575737 358400
rect 575771 358366 575777 358400
rect 575731 358328 575777 358366
rect 575731 358294 575737 358328
rect 575771 358294 575777 358328
rect 575731 358256 575777 358294
rect 575731 358222 575737 358256
rect 575771 358222 575777 358256
rect 575731 358184 575777 358222
rect 575731 358150 575737 358184
rect 575771 358150 575777 358184
rect 575731 358112 575777 358150
rect 575731 358078 575737 358112
rect 575771 358078 575777 358112
rect 575731 358040 575777 358078
rect 575731 358006 575737 358040
rect 575771 358006 575777 358040
rect 575731 357968 575777 358006
rect 575731 357934 575737 357968
rect 575771 357934 575777 357968
rect 575731 357919 575777 357934
rect 575989 358904 576035 358919
rect 575989 358870 575995 358904
rect 576029 358870 576035 358904
rect 575989 358832 576035 358870
rect 575989 358798 575995 358832
rect 576029 358798 576035 358832
rect 575989 358760 576035 358798
rect 575989 358726 575995 358760
rect 576029 358726 576035 358760
rect 575989 358688 576035 358726
rect 575989 358654 575995 358688
rect 576029 358654 576035 358688
rect 575989 358616 576035 358654
rect 575989 358582 575995 358616
rect 576029 358582 576035 358616
rect 575989 358544 576035 358582
rect 575989 358510 575995 358544
rect 576029 358510 576035 358544
rect 575989 358472 576035 358510
rect 575989 358438 575995 358472
rect 576029 358438 576035 358472
rect 575989 358400 576035 358438
rect 575989 358366 575995 358400
rect 576029 358366 576035 358400
rect 575989 358328 576035 358366
rect 575989 358294 575995 358328
rect 576029 358294 576035 358328
rect 575989 358256 576035 358294
rect 575989 358222 575995 358256
rect 576029 358222 576035 358256
rect 575989 358184 576035 358222
rect 575989 358150 575995 358184
rect 576029 358150 576035 358184
rect 575989 358112 576035 358150
rect 575989 358078 575995 358112
rect 576029 358078 576035 358112
rect 575989 358040 576035 358078
rect 575989 358006 575995 358040
rect 576029 358006 576035 358040
rect 575989 357968 576035 358006
rect 575989 357934 575995 357968
rect 576029 357934 576035 357968
rect 575989 357919 576035 357934
rect 576247 358904 576293 358919
rect 576247 358870 576253 358904
rect 576287 358870 576293 358904
rect 576247 358832 576293 358870
rect 576247 358798 576253 358832
rect 576287 358798 576293 358832
rect 576247 358760 576293 358798
rect 576247 358726 576253 358760
rect 576287 358726 576293 358760
rect 576247 358688 576293 358726
rect 576247 358654 576253 358688
rect 576287 358654 576293 358688
rect 576247 358616 576293 358654
rect 576247 358582 576253 358616
rect 576287 358582 576293 358616
rect 576247 358544 576293 358582
rect 576247 358510 576253 358544
rect 576287 358510 576293 358544
rect 576247 358472 576293 358510
rect 576247 358438 576253 358472
rect 576287 358438 576293 358472
rect 576247 358400 576293 358438
rect 576247 358366 576253 358400
rect 576287 358366 576293 358400
rect 576247 358328 576293 358366
rect 576247 358294 576253 358328
rect 576287 358294 576293 358328
rect 576247 358256 576293 358294
rect 576247 358222 576253 358256
rect 576287 358222 576293 358256
rect 576247 358184 576293 358222
rect 576247 358150 576253 358184
rect 576287 358150 576293 358184
rect 576247 358112 576293 358150
rect 576247 358078 576253 358112
rect 576287 358078 576293 358112
rect 576247 358040 576293 358078
rect 576247 358006 576253 358040
rect 576287 358006 576293 358040
rect 576247 357968 576293 358006
rect 576247 357934 576253 357968
rect 576287 357934 576293 357968
rect 576247 357919 576293 357934
rect 576505 358904 576551 358919
rect 576505 358870 576511 358904
rect 576545 358870 576551 358904
rect 576505 358832 576551 358870
rect 576505 358798 576511 358832
rect 576545 358798 576551 358832
rect 576505 358760 576551 358798
rect 576505 358726 576511 358760
rect 576545 358726 576551 358760
rect 576505 358688 576551 358726
rect 576505 358654 576511 358688
rect 576545 358654 576551 358688
rect 576505 358616 576551 358654
rect 576505 358582 576511 358616
rect 576545 358582 576551 358616
rect 576505 358544 576551 358582
rect 576505 358510 576511 358544
rect 576545 358510 576551 358544
rect 576505 358472 576551 358510
rect 576505 358438 576511 358472
rect 576545 358438 576551 358472
rect 576505 358400 576551 358438
rect 576505 358366 576511 358400
rect 576545 358366 576551 358400
rect 576505 358328 576551 358366
rect 576505 358294 576511 358328
rect 576545 358294 576551 358328
rect 576505 358256 576551 358294
rect 576505 358222 576511 358256
rect 576545 358222 576551 358256
rect 576505 358184 576551 358222
rect 576505 358150 576511 358184
rect 576545 358150 576551 358184
rect 576505 358112 576551 358150
rect 576505 358078 576511 358112
rect 576545 358078 576551 358112
rect 576505 358040 576551 358078
rect 576505 358006 576511 358040
rect 576545 358006 576551 358040
rect 576505 357968 576551 358006
rect 576505 357934 576511 357968
rect 576545 357934 576551 357968
rect 576505 357919 576551 357934
rect 576763 358904 576809 358919
rect 576763 358870 576769 358904
rect 576803 358870 576809 358904
rect 576763 358832 576809 358870
rect 576763 358798 576769 358832
rect 576803 358798 576809 358832
rect 576763 358760 576809 358798
rect 576763 358726 576769 358760
rect 576803 358726 576809 358760
rect 576763 358688 576809 358726
rect 576763 358654 576769 358688
rect 576803 358654 576809 358688
rect 576763 358616 576809 358654
rect 576763 358582 576769 358616
rect 576803 358582 576809 358616
rect 576763 358544 576809 358582
rect 576763 358510 576769 358544
rect 576803 358510 576809 358544
rect 576763 358472 576809 358510
rect 576763 358438 576769 358472
rect 576803 358438 576809 358472
rect 576763 358400 576809 358438
rect 576763 358366 576769 358400
rect 576803 358366 576809 358400
rect 576763 358328 576809 358366
rect 576763 358294 576769 358328
rect 576803 358294 576809 358328
rect 576763 358256 576809 358294
rect 576763 358222 576769 358256
rect 576803 358222 576809 358256
rect 576763 358184 576809 358222
rect 576763 358150 576769 358184
rect 576803 358150 576809 358184
rect 576763 358112 576809 358150
rect 576763 358078 576769 358112
rect 576803 358078 576809 358112
rect 576763 358040 576809 358078
rect 576763 358006 576769 358040
rect 576803 358006 576809 358040
rect 576763 357968 576809 358006
rect 576763 357934 576769 357968
rect 576803 357934 576809 357968
rect 576763 357919 576809 357934
rect 577021 358904 577067 358919
rect 577021 358870 577027 358904
rect 577061 358870 577067 358904
rect 577021 358832 577067 358870
rect 577021 358798 577027 358832
rect 577061 358798 577067 358832
rect 577021 358760 577067 358798
rect 577021 358726 577027 358760
rect 577061 358726 577067 358760
rect 577021 358688 577067 358726
rect 577021 358654 577027 358688
rect 577061 358654 577067 358688
rect 577021 358616 577067 358654
rect 577021 358582 577027 358616
rect 577061 358582 577067 358616
rect 577021 358544 577067 358582
rect 577021 358510 577027 358544
rect 577061 358510 577067 358544
rect 577021 358472 577067 358510
rect 577021 358438 577027 358472
rect 577061 358438 577067 358472
rect 577021 358400 577067 358438
rect 577021 358366 577027 358400
rect 577061 358366 577067 358400
rect 577021 358328 577067 358366
rect 577021 358294 577027 358328
rect 577061 358294 577067 358328
rect 577021 358256 577067 358294
rect 577021 358222 577027 358256
rect 577061 358222 577067 358256
rect 577021 358184 577067 358222
rect 577021 358150 577027 358184
rect 577061 358150 577067 358184
rect 577021 358112 577067 358150
rect 577021 358078 577027 358112
rect 577061 358078 577067 358112
rect 577021 358040 577067 358078
rect 577021 358006 577027 358040
rect 577061 358006 577067 358040
rect 577021 357968 577067 358006
rect 577021 357934 577027 357968
rect 577061 357934 577067 357968
rect 577021 357919 577067 357934
rect 577279 358904 577325 358919
rect 577279 358870 577285 358904
rect 577319 358870 577325 358904
rect 577279 358832 577325 358870
rect 577279 358798 577285 358832
rect 577319 358798 577325 358832
rect 577279 358760 577325 358798
rect 577279 358726 577285 358760
rect 577319 358726 577325 358760
rect 577279 358688 577325 358726
rect 577279 358654 577285 358688
rect 577319 358654 577325 358688
rect 577279 358616 577325 358654
rect 577279 358582 577285 358616
rect 577319 358582 577325 358616
rect 577279 358544 577325 358582
rect 577279 358510 577285 358544
rect 577319 358510 577325 358544
rect 577279 358472 577325 358510
rect 577279 358438 577285 358472
rect 577319 358438 577325 358472
rect 577279 358400 577325 358438
rect 577279 358366 577285 358400
rect 577319 358366 577325 358400
rect 577279 358328 577325 358366
rect 577279 358294 577285 358328
rect 577319 358294 577325 358328
rect 577279 358256 577325 358294
rect 577279 358222 577285 358256
rect 577319 358222 577325 358256
rect 577279 358184 577325 358222
rect 577279 358150 577285 358184
rect 577319 358150 577325 358184
rect 577279 358112 577325 358150
rect 577279 358078 577285 358112
rect 577319 358078 577325 358112
rect 577279 358040 577325 358078
rect 577279 358006 577285 358040
rect 577319 358006 577325 358040
rect 577279 357968 577325 358006
rect 577279 357934 577285 357968
rect 577319 357934 577325 357968
rect 577279 357919 577325 357934
rect 577537 358904 577583 358919
rect 577537 358870 577543 358904
rect 577577 358870 577583 358904
rect 577537 358832 577583 358870
rect 577537 358798 577543 358832
rect 577577 358798 577583 358832
rect 577537 358760 577583 358798
rect 577537 358726 577543 358760
rect 577577 358726 577583 358760
rect 577537 358688 577583 358726
rect 577537 358654 577543 358688
rect 577577 358654 577583 358688
rect 577537 358616 577583 358654
rect 577537 358582 577543 358616
rect 577577 358582 577583 358616
rect 577537 358544 577583 358582
rect 577537 358510 577543 358544
rect 577577 358510 577583 358544
rect 577537 358472 577583 358510
rect 577537 358438 577543 358472
rect 577577 358438 577583 358472
rect 577537 358400 577583 358438
rect 577537 358366 577543 358400
rect 577577 358366 577583 358400
rect 577537 358328 577583 358366
rect 577537 358294 577543 358328
rect 577577 358294 577583 358328
rect 577537 358256 577583 358294
rect 577537 358222 577543 358256
rect 577577 358222 577583 358256
rect 577537 358184 577583 358222
rect 577537 358150 577543 358184
rect 577577 358150 577583 358184
rect 577537 358112 577583 358150
rect 577537 358078 577543 358112
rect 577577 358078 577583 358112
rect 577537 358040 577583 358078
rect 577537 358006 577543 358040
rect 577577 358006 577583 358040
rect 577537 357968 577583 358006
rect 577537 357934 577543 357968
rect 577577 357934 577583 357968
rect 577537 357919 577583 357934
rect 577795 358904 577841 358919
rect 577795 358870 577801 358904
rect 577835 358870 577841 358904
rect 577795 358832 577841 358870
rect 577795 358798 577801 358832
rect 577835 358798 577841 358832
rect 577795 358760 577841 358798
rect 577795 358726 577801 358760
rect 577835 358726 577841 358760
rect 577795 358688 577841 358726
rect 577795 358654 577801 358688
rect 577835 358654 577841 358688
rect 577795 358616 577841 358654
rect 577795 358582 577801 358616
rect 577835 358582 577841 358616
rect 577795 358544 577841 358582
rect 577795 358510 577801 358544
rect 577835 358510 577841 358544
rect 577795 358472 577841 358510
rect 577795 358438 577801 358472
rect 577835 358438 577841 358472
rect 577795 358400 577841 358438
rect 577795 358366 577801 358400
rect 577835 358366 577841 358400
rect 577795 358328 577841 358366
rect 577795 358294 577801 358328
rect 577835 358294 577841 358328
rect 577795 358256 577841 358294
rect 577795 358222 577801 358256
rect 577835 358222 577841 358256
rect 577795 358184 577841 358222
rect 577795 358150 577801 358184
rect 577835 358150 577841 358184
rect 577795 358112 577841 358150
rect 577795 358078 577801 358112
rect 577835 358078 577841 358112
rect 577795 358040 577841 358078
rect 577795 358006 577801 358040
rect 577835 358006 577841 358040
rect 577795 357968 577841 358006
rect 577795 357934 577801 357968
rect 577835 357934 577841 357968
rect 577795 357919 577841 357934
rect 578053 358904 578099 358919
rect 578053 358870 578059 358904
rect 578093 358870 578099 358904
rect 578053 358832 578099 358870
rect 578053 358798 578059 358832
rect 578093 358798 578099 358832
rect 578053 358760 578099 358798
rect 578053 358726 578059 358760
rect 578093 358726 578099 358760
rect 578053 358688 578099 358726
rect 578053 358654 578059 358688
rect 578093 358654 578099 358688
rect 578053 358616 578099 358654
rect 578053 358582 578059 358616
rect 578093 358582 578099 358616
rect 578053 358544 578099 358582
rect 578053 358510 578059 358544
rect 578093 358510 578099 358544
rect 578053 358472 578099 358510
rect 578053 358438 578059 358472
rect 578093 358438 578099 358472
rect 578053 358400 578099 358438
rect 578053 358366 578059 358400
rect 578093 358366 578099 358400
rect 578053 358328 578099 358366
rect 578053 358294 578059 358328
rect 578093 358294 578099 358328
rect 578053 358256 578099 358294
rect 578053 358222 578059 358256
rect 578093 358222 578099 358256
rect 578053 358184 578099 358222
rect 578053 358150 578059 358184
rect 578093 358150 578099 358184
rect 578053 358112 578099 358150
rect 578053 358078 578059 358112
rect 578093 358078 578099 358112
rect 578053 358040 578099 358078
rect 578053 358006 578059 358040
rect 578093 358006 578099 358040
rect 578053 357968 578099 358006
rect 578053 357934 578059 357968
rect 578093 357934 578099 357968
rect 578053 357919 578099 357934
rect 578311 358904 578357 358919
rect 578311 358870 578317 358904
rect 578351 358870 578357 358904
rect 578311 358832 578357 358870
rect 578311 358798 578317 358832
rect 578351 358798 578357 358832
rect 578311 358760 578357 358798
rect 578311 358726 578317 358760
rect 578351 358726 578357 358760
rect 578311 358688 578357 358726
rect 578311 358654 578317 358688
rect 578351 358654 578357 358688
rect 578311 358616 578357 358654
rect 578311 358582 578317 358616
rect 578351 358582 578357 358616
rect 578311 358544 578357 358582
rect 578311 358510 578317 358544
rect 578351 358510 578357 358544
rect 578311 358472 578357 358510
rect 578311 358438 578317 358472
rect 578351 358438 578357 358472
rect 578311 358400 578357 358438
rect 578311 358366 578317 358400
rect 578351 358366 578357 358400
rect 578311 358328 578357 358366
rect 578311 358294 578317 358328
rect 578351 358294 578357 358328
rect 578311 358256 578357 358294
rect 578311 358222 578317 358256
rect 578351 358222 578357 358256
rect 578311 358184 578357 358222
rect 578311 358150 578317 358184
rect 578351 358150 578357 358184
rect 578311 358112 578357 358150
rect 578311 358078 578317 358112
rect 578351 358078 578357 358112
rect 578311 358040 578357 358078
rect 578311 358006 578317 358040
rect 578351 358006 578357 358040
rect 578311 357968 578357 358006
rect 578311 357934 578317 357968
rect 578351 357934 578357 357968
rect 578311 357919 578357 357934
rect 578569 358904 578615 358919
rect 578569 358870 578575 358904
rect 578609 358870 578615 358904
rect 578569 358832 578615 358870
rect 578569 358798 578575 358832
rect 578609 358798 578615 358832
rect 578569 358760 578615 358798
rect 578569 358726 578575 358760
rect 578609 358726 578615 358760
rect 578569 358688 578615 358726
rect 578569 358654 578575 358688
rect 578609 358654 578615 358688
rect 578569 358616 578615 358654
rect 578569 358582 578575 358616
rect 578609 358582 578615 358616
rect 578569 358544 578615 358582
rect 578569 358510 578575 358544
rect 578609 358510 578615 358544
rect 578569 358472 578615 358510
rect 578569 358438 578575 358472
rect 578609 358438 578615 358472
rect 578569 358400 578615 358438
rect 578569 358366 578575 358400
rect 578609 358366 578615 358400
rect 578569 358328 578615 358366
rect 578569 358294 578575 358328
rect 578609 358294 578615 358328
rect 578569 358256 578615 358294
rect 578569 358222 578575 358256
rect 578609 358222 578615 358256
rect 578569 358184 578615 358222
rect 578569 358150 578575 358184
rect 578609 358150 578615 358184
rect 578569 358112 578615 358150
rect 578569 358078 578575 358112
rect 578609 358078 578615 358112
rect 578569 358040 578615 358078
rect 578569 358006 578575 358040
rect 578609 358006 578615 358040
rect 578569 357968 578615 358006
rect 578569 357934 578575 357968
rect 578609 357934 578615 357968
rect 578569 357919 578615 357934
rect 578827 358904 578873 358919
rect 578827 358870 578833 358904
rect 578867 358870 578873 358904
rect 578827 358832 578873 358870
rect 578827 358798 578833 358832
rect 578867 358798 578873 358832
rect 578827 358760 578873 358798
rect 578827 358726 578833 358760
rect 578867 358726 578873 358760
rect 578827 358688 578873 358726
rect 578827 358654 578833 358688
rect 578867 358654 578873 358688
rect 578827 358616 578873 358654
rect 578827 358582 578833 358616
rect 578867 358582 578873 358616
rect 578827 358544 578873 358582
rect 578827 358510 578833 358544
rect 578867 358510 578873 358544
rect 578827 358472 578873 358510
rect 578827 358438 578833 358472
rect 578867 358438 578873 358472
rect 578827 358400 578873 358438
rect 578827 358366 578833 358400
rect 578867 358366 578873 358400
rect 578827 358328 578873 358366
rect 578827 358294 578833 358328
rect 578867 358294 578873 358328
rect 578827 358256 578873 358294
rect 578827 358222 578833 358256
rect 578867 358222 578873 358256
rect 578827 358184 578873 358222
rect 578827 358150 578833 358184
rect 578867 358150 578873 358184
rect 578827 358112 578873 358150
rect 578827 358078 578833 358112
rect 578867 358078 578873 358112
rect 578827 358040 578873 358078
rect 578827 358006 578833 358040
rect 578867 358006 578873 358040
rect 578827 357968 578873 358006
rect 578827 357934 578833 357968
rect 578867 357934 578873 357968
rect 578827 357919 578873 357934
rect 579085 358904 579131 358919
rect 579085 358870 579091 358904
rect 579125 358870 579131 358904
rect 579085 358832 579131 358870
rect 579085 358798 579091 358832
rect 579125 358798 579131 358832
rect 579085 358760 579131 358798
rect 579085 358726 579091 358760
rect 579125 358726 579131 358760
rect 579085 358688 579131 358726
rect 579085 358654 579091 358688
rect 579125 358654 579131 358688
rect 579085 358616 579131 358654
rect 579085 358582 579091 358616
rect 579125 358582 579131 358616
rect 579085 358544 579131 358582
rect 579085 358510 579091 358544
rect 579125 358510 579131 358544
rect 579085 358472 579131 358510
rect 579085 358438 579091 358472
rect 579125 358438 579131 358472
rect 579085 358400 579131 358438
rect 579085 358366 579091 358400
rect 579125 358366 579131 358400
rect 579085 358328 579131 358366
rect 579085 358294 579091 358328
rect 579125 358294 579131 358328
rect 579085 358256 579131 358294
rect 579085 358222 579091 358256
rect 579125 358222 579131 358256
rect 579085 358184 579131 358222
rect 579085 358150 579091 358184
rect 579125 358150 579131 358184
rect 579085 358112 579131 358150
rect 579085 358078 579091 358112
rect 579125 358078 579131 358112
rect 579085 358040 579131 358078
rect 579085 358006 579091 358040
rect 579125 358006 579131 358040
rect 579085 357968 579131 358006
rect 579085 357934 579091 357968
rect 579125 357934 579131 357968
rect 579085 357919 579131 357934
rect 579343 358904 579389 358919
rect 579343 358870 579349 358904
rect 579383 358870 579389 358904
rect 579343 358832 579389 358870
rect 579343 358798 579349 358832
rect 579383 358798 579389 358832
rect 579343 358760 579389 358798
rect 579343 358726 579349 358760
rect 579383 358726 579389 358760
rect 579343 358688 579389 358726
rect 579343 358654 579349 358688
rect 579383 358654 579389 358688
rect 579343 358616 579389 358654
rect 579343 358582 579349 358616
rect 579383 358582 579389 358616
rect 579343 358544 579389 358582
rect 579343 358510 579349 358544
rect 579383 358510 579389 358544
rect 579343 358472 579389 358510
rect 579343 358438 579349 358472
rect 579383 358438 579389 358472
rect 579343 358400 579389 358438
rect 579343 358366 579349 358400
rect 579383 358366 579389 358400
rect 579343 358328 579389 358366
rect 579343 358294 579349 358328
rect 579383 358294 579389 358328
rect 579343 358256 579389 358294
rect 579343 358222 579349 358256
rect 579383 358222 579389 358256
rect 579343 358184 579389 358222
rect 579343 358150 579349 358184
rect 579383 358150 579389 358184
rect 579343 358112 579389 358150
rect 579343 358078 579349 358112
rect 579383 358078 579389 358112
rect 579343 358040 579389 358078
rect 579343 358006 579349 358040
rect 579383 358006 579389 358040
rect 579343 357968 579389 358006
rect 579343 357934 579349 357968
rect 579383 357934 579389 357968
rect 579343 357919 579389 357934
rect 579601 358904 579647 358919
rect 579601 358870 579607 358904
rect 579641 358870 579647 358904
rect 579601 358832 579647 358870
rect 579601 358798 579607 358832
rect 579641 358798 579647 358832
rect 579601 358760 579647 358798
rect 579601 358726 579607 358760
rect 579641 358726 579647 358760
rect 579601 358688 579647 358726
rect 579601 358654 579607 358688
rect 579641 358654 579647 358688
rect 579601 358616 579647 358654
rect 579601 358582 579607 358616
rect 579641 358582 579647 358616
rect 579601 358544 579647 358582
rect 579601 358510 579607 358544
rect 579641 358510 579647 358544
rect 579601 358472 579647 358510
rect 579601 358438 579607 358472
rect 579641 358438 579647 358472
rect 579601 358400 579647 358438
rect 579601 358366 579607 358400
rect 579641 358366 579647 358400
rect 579601 358328 579647 358366
rect 579601 358294 579607 358328
rect 579641 358294 579647 358328
rect 579601 358256 579647 358294
rect 579601 358222 579607 358256
rect 579641 358222 579647 358256
rect 579601 358184 579647 358222
rect 579601 358150 579607 358184
rect 579641 358150 579647 358184
rect 579601 358112 579647 358150
rect 579601 358078 579607 358112
rect 579641 358078 579647 358112
rect 579601 358040 579647 358078
rect 579601 358006 579607 358040
rect 579641 358006 579647 358040
rect 579601 357968 579647 358006
rect 579601 357934 579607 357968
rect 579641 357934 579647 357968
rect 579601 357919 579647 357934
rect 579859 358904 579905 358919
rect 579859 358870 579865 358904
rect 579899 358870 579905 358904
rect 579859 358832 579905 358870
rect 579859 358798 579865 358832
rect 579899 358798 579905 358832
rect 579859 358760 579905 358798
rect 579859 358726 579865 358760
rect 579899 358726 579905 358760
rect 579859 358688 579905 358726
rect 579859 358654 579865 358688
rect 579899 358654 579905 358688
rect 579859 358616 579905 358654
rect 579859 358582 579865 358616
rect 579899 358582 579905 358616
rect 579859 358544 579905 358582
rect 579859 358510 579865 358544
rect 579899 358510 579905 358544
rect 579859 358472 579905 358510
rect 579859 358438 579865 358472
rect 579899 358438 579905 358472
rect 579859 358400 579905 358438
rect 579859 358366 579865 358400
rect 579899 358366 579905 358400
rect 579859 358328 579905 358366
rect 579859 358294 579865 358328
rect 579899 358294 579905 358328
rect 579859 358256 579905 358294
rect 579859 358222 579865 358256
rect 579899 358222 579905 358256
rect 579859 358184 579905 358222
rect 579859 358150 579865 358184
rect 579899 358150 579905 358184
rect 579859 358112 579905 358150
rect 579859 358078 579865 358112
rect 579899 358078 579905 358112
rect 579859 358040 579905 358078
rect 579859 358006 579865 358040
rect 579899 358006 579905 358040
rect 579859 357968 579905 358006
rect 579859 357934 579865 357968
rect 579899 357934 579905 357968
rect 579859 357919 579905 357934
rect 580266 357835 580370 359795
rect 573877 357691 574526 357819
rect 580018 357796 580370 357835
rect 580018 357762 580058 357796
rect 580092 357762 580370 357796
rect 580018 357731 580370 357762
rect 580018 357729 580132 357731
rect 573877 357654 574522 357691
rect 573877 357620 574451 357654
rect 574485 357620 574522 357654
rect 573877 357612 574522 357620
rect 573523 357573 574522 357612
rect 565774 357549 566084 357551
rect 559746 357506 566084 357549
rect 559746 357472 560755 357506
rect 560789 357472 560955 357506
rect 560989 357472 561155 357506
rect 561189 357472 561355 357506
rect 561389 357472 561555 357506
rect 561589 357472 561755 357506
rect 561789 357472 561955 357506
rect 561989 357472 562155 357506
rect 562189 357472 562355 357506
rect 562389 357472 562555 357506
rect 562589 357472 562755 357506
rect 562789 357472 562955 357506
rect 562989 357472 563155 357506
rect 563189 357472 563355 357506
rect 563389 357472 563555 357506
rect 563589 357472 563755 357506
rect 563789 357472 563955 357506
rect 563989 357472 564155 357506
rect 564189 357472 564355 357506
rect 564389 357472 564555 357506
rect 564589 357472 564755 357506
rect 564789 357472 564955 357506
rect 564989 357472 565155 357506
rect 565189 357472 565355 357506
rect 565389 357472 565555 357506
rect 565589 357472 566084 357506
rect 559746 357431 566084 357472
rect 559746 357429 565870 357431
rect 565964 357239 566084 357431
rect 574658 357436 580044 357479
rect 574658 357402 574729 357436
rect 574763 357402 574929 357436
rect 574963 357402 575129 357436
rect 575163 357402 575329 357436
rect 575363 357402 575529 357436
rect 575563 357402 575729 357436
rect 575763 357402 575929 357436
rect 575963 357402 576129 357436
rect 576163 357402 576329 357436
rect 576363 357402 576529 357436
rect 576563 357402 576729 357436
rect 576763 357402 576929 357436
rect 576963 357402 577129 357436
rect 577163 357402 577329 357436
rect 577363 357402 577529 357436
rect 577563 357402 577729 357436
rect 577763 357402 577929 357436
rect 577963 357402 578129 357436
rect 578163 357402 578329 357436
rect 578363 357402 578529 357436
rect 578563 357402 578729 357436
rect 578763 357402 578929 357436
rect 578963 357402 579129 357436
rect 579163 357402 579329 357436
rect 579363 357402 579529 357436
rect 579563 357402 579729 357436
rect 579763 357402 580044 357436
rect 574658 357359 580044 357402
rect 574776 357239 574896 357359
rect 565964 357119 574896 357239
rect 508600 356609 508756 356611
rect 508600 356429 508620 356609
rect 508736 356429 508756 356609
rect 508600 356427 508756 356429
rect 565612 314307 573784 314427
rect 565612 313121 565732 314307
rect 560418 313078 565732 313121
rect 560418 313044 560617 313078
rect 560651 313044 560817 313078
rect 560851 313044 561017 313078
rect 561051 313044 561217 313078
rect 561251 313044 561417 313078
rect 561451 313044 561617 313078
rect 561651 313044 561817 313078
rect 561851 313044 562017 313078
rect 562051 313044 562217 313078
rect 562251 313044 562417 313078
rect 562451 313044 562617 313078
rect 562651 313044 562817 313078
rect 562851 313044 563017 313078
rect 563051 313044 563217 313078
rect 563251 313044 563417 313078
rect 563451 313044 563617 313078
rect 563651 313044 563817 313078
rect 563851 313044 564017 313078
rect 564051 313044 564217 313078
rect 564251 313044 564417 313078
rect 564451 313044 564617 313078
rect 564651 313044 564817 313078
rect 564851 313044 565017 313078
rect 565051 313044 565217 313078
rect 565251 313044 565417 313078
rect 565451 313044 565732 313078
rect 560418 313001 565732 313044
rect 566130 313806 566370 313813
rect 566130 313626 566160 313806
rect 566340 313803 566370 313806
rect 566340 313626 566376 313803
rect 560423 312666 560469 312681
rect 560423 312632 560429 312666
rect 560463 312632 560469 312666
rect 560423 312594 560469 312632
rect 560423 312560 560429 312594
rect 560463 312560 560469 312594
rect 560423 312522 560469 312560
rect 560423 312488 560429 312522
rect 560463 312488 560469 312522
rect 560423 312450 560469 312488
rect 560423 312416 560429 312450
rect 560463 312416 560469 312450
rect 560423 312378 560469 312416
rect 560423 312344 560429 312378
rect 560463 312344 560469 312378
rect 560423 312306 560469 312344
rect 560423 312272 560429 312306
rect 560463 312272 560469 312306
rect 560423 312234 560469 312272
rect 560423 312200 560429 312234
rect 560463 312200 560469 312234
rect 560423 312162 560469 312200
rect 560423 312128 560429 312162
rect 560463 312128 560469 312162
rect 560423 312090 560469 312128
rect 560423 312056 560429 312090
rect 560463 312056 560469 312090
rect 560423 312018 560469 312056
rect 560423 311984 560429 312018
rect 560463 311984 560469 312018
rect 560423 311946 560469 311984
rect 560423 311912 560429 311946
rect 560463 311912 560469 311946
rect 560423 311874 560469 311912
rect 560423 311840 560429 311874
rect 560463 311840 560469 311874
rect 560423 311802 560469 311840
rect 560423 311768 560429 311802
rect 560463 311768 560469 311802
rect 559656 311739 560254 311753
rect 559656 311559 559680 311739
rect 559860 311701 560254 311739
rect 559860 311595 560121 311701
rect 560227 311595 560254 311701
rect 560423 311730 560469 311768
rect 560423 311696 560429 311730
rect 560463 311696 560469 311730
rect 560423 311681 560469 311696
rect 560681 312666 560727 312681
rect 560681 312632 560687 312666
rect 560721 312632 560727 312666
rect 560681 312594 560727 312632
rect 560681 312560 560687 312594
rect 560721 312560 560727 312594
rect 560681 312522 560727 312560
rect 560681 312488 560687 312522
rect 560721 312488 560727 312522
rect 560681 312450 560727 312488
rect 560681 312416 560687 312450
rect 560721 312416 560727 312450
rect 560681 312378 560727 312416
rect 560681 312344 560687 312378
rect 560721 312344 560727 312378
rect 560681 312306 560727 312344
rect 560681 312272 560687 312306
rect 560721 312272 560727 312306
rect 560681 312234 560727 312272
rect 560681 312200 560687 312234
rect 560721 312200 560727 312234
rect 560681 312162 560727 312200
rect 560681 312128 560687 312162
rect 560721 312128 560727 312162
rect 560681 312090 560727 312128
rect 560681 312056 560687 312090
rect 560721 312056 560727 312090
rect 560681 312018 560727 312056
rect 560681 311984 560687 312018
rect 560721 311984 560727 312018
rect 560681 311946 560727 311984
rect 560681 311912 560687 311946
rect 560721 311912 560727 311946
rect 560681 311874 560727 311912
rect 560681 311840 560687 311874
rect 560721 311840 560727 311874
rect 560681 311802 560727 311840
rect 560681 311768 560687 311802
rect 560721 311768 560727 311802
rect 560681 311730 560727 311768
rect 560681 311696 560687 311730
rect 560721 311696 560727 311730
rect 560681 311681 560727 311696
rect 560939 312666 560985 312681
rect 560939 312632 560945 312666
rect 560979 312632 560985 312666
rect 560939 312594 560985 312632
rect 560939 312560 560945 312594
rect 560979 312560 560985 312594
rect 560939 312522 560985 312560
rect 560939 312488 560945 312522
rect 560979 312488 560985 312522
rect 560939 312450 560985 312488
rect 560939 312416 560945 312450
rect 560979 312416 560985 312450
rect 560939 312378 560985 312416
rect 560939 312344 560945 312378
rect 560979 312344 560985 312378
rect 560939 312306 560985 312344
rect 560939 312272 560945 312306
rect 560979 312272 560985 312306
rect 560939 312234 560985 312272
rect 560939 312200 560945 312234
rect 560979 312200 560985 312234
rect 560939 312162 560985 312200
rect 560939 312128 560945 312162
rect 560979 312128 560985 312162
rect 560939 312090 560985 312128
rect 560939 312056 560945 312090
rect 560979 312056 560985 312090
rect 560939 312018 560985 312056
rect 560939 311984 560945 312018
rect 560979 311984 560985 312018
rect 560939 311946 560985 311984
rect 560939 311912 560945 311946
rect 560979 311912 560985 311946
rect 560939 311874 560985 311912
rect 560939 311840 560945 311874
rect 560979 311840 560985 311874
rect 560939 311802 560985 311840
rect 560939 311768 560945 311802
rect 560979 311768 560985 311802
rect 560939 311730 560985 311768
rect 560939 311696 560945 311730
rect 560979 311696 560985 311730
rect 560939 311681 560985 311696
rect 561197 312666 561243 312681
rect 561197 312632 561203 312666
rect 561237 312632 561243 312666
rect 561197 312594 561243 312632
rect 561197 312560 561203 312594
rect 561237 312560 561243 312594
rect 561197 312522 561243 312560
rect 561197 312488 561203 312522
rect 561237 312488 561243 312522
rect 561197 312450 561243 312488
rect 561197 312416 561203 312450
rect 561237 312416 561243 312450
rect 561197 312378 561243 312416
rect 561197 312344 561203 312378
rect 561237 312344 561243 312378
rect 561197 312306 561243 312344
rect 561197 312272 561203 312306
rect 561237 312272 561243 312306
rect 561197 312234 561243 312272
rect 561197 312200 561203 312234
rect 561237 312200 561243 312234
rect 561197 312162 561243 312200
rect 561197 312128 561203 312162
rect 561237 312128 561243 312162
rect 561197 312090 561243 312128
rect 561197 312056 561203 312090
rect 561237 312056 561243 312090
rect 561197 312018 561243 312056
rect 561197 311984 561203 312018
rect 561237 311984 561243 312018
rect 561197 311946 561243 311984
rect 561197 311912 561203 311946
rect 561237 311912 561243 311946
rect 561197 311874 561243 311912
rect 561197 311840 561203 311874
rect 561237 311840 561243 311874
rect 561197 311802 561243 311840
rect 561197 311768 561203 311802
rect 561237 311768 561243 311802
rect 561197 311730 561243 311768
rect 561197 311696 561203 311730
rect 561237 311696 561243 311730
rect 561197 311681 561243 311696
rect 561455 312666 561501 312681
rect 561455 312632 561461 312666
rect 561495 312632 561501 312666
rect 561455 312594 561501 312632
rect 561455 312560 561461 312594
rect 561495 312560 561501 312594
rect 561455 312522 561501 312560
rect 561455 312488 561461 312522
rect 561495 312488 561501 312522
rect 561455 312450 561501 312488
rect 561455 312416 561461 312450
rect 561495 312416 561501 312450
rect 561455 312378 561501 312416
rect 561455 312344 561461 312378
rect 561495 312344 561501 312378
rect 561455 312306 561501 312344
rect 561455 312272 561461 312306
rect 561495 312272 561501 312306
rect 561455 312234 561501 312272
rect 561455 312200 561461 312234
rect 561495 312200 561501 312234
rect 561455 312162 561501 312200
rect 561455 312128 561461 312162
rect 561495 312128 561501 312162
rect 561455 312090 561501 312128
rect 561455 312056 561461 312090
rect 561495 312056 561501 312090
rect 561455 312018 561501 312056
rect 561455 311984 561461 312018
rect 561495 311984 561501 312018
rect 561455 311946 561501 311984
rect 561455 311912 561461 311946
rect 561495 311912 561501 311946
rect 561455 311874 561501 311912
rect 561455 311840 561461 311874
rect 561495 311840 561501 311874
rect 561455 311802 561501 311840
rect 561455 311768 561461 311802
rect 561495 311768 561501 311802
rect 561455 311730 561501 311768
rect 561455 311696 561461 311730
rect 561495 311696 561501 311730
rect 561455 311681 561501 311696
rect 561713 312666 561759 312681
rect 561713 312632 561719 312666
rect 561753 312632 561759 312666
rect 561713 312594 561759 312632
rect 561713 312560 561719 312594
rect 561753 312560 561759 312594
rect 561713 312522 561759 312560
rect 561713 312488 561719 312522
rect 561753 312488 561759 312522
rect 561713 312450 561759 312488
rect 561713 312416 561719 312450
rect 561753 312416 561759 312450
rect 561713 312378 561759 312416
rect 561713 312344 561719 312378
rect 561753 312344 561759 312378
rect 561713 312306 561759 312344
rect 561713 312272 561719 312306
rect 561753 312272 561759 312306
rect 561713 312234 561759 312272
rect 561713 312200 561719 312234
rect 561753 312200 561759 312234
rect 561713 312162 561759 312200
rect 561713 312128 561719 312162
rect 561753 312128 561759 312162
rect 561713 312090 561759 312128
rect 561713 312056 561719 312090
rect 561753 312056 561759 312090
rect 561713 312018 561759 312056
rect 561713 311984 561719 312018
rect 561753 311984 561759 312018
rect 561713 311946 561759 311984
rect 561713 311912 561719 311946
rect 561753 311912 561759 311946
rect 561713 311874 561759 311912
rect 561713 311840 561719 311874
rect 561753 311840 561759 311874
rect 561713 311802 561759 311840
rect 561713 311768 561719 311802
rect 561753 311768 561759 311802
rect 561713 311730 561759 311768
rect 561713 311696 561719 311730
rect 561753 311696 561759 311730
rect 561713 311681 561759 311696
rect 561971 312666 562017 312681
rect 561971 312632 561977 312666
rect 562011 312632 562017 312666
rect 561971 312594 562017 312632
rect 561971 312560 561977 312594
rect 562011 312560 562017 312594
rect 561971 312522 562017 312560
rect 561971 312488 561977 312522
rect 562011 312488 562017 312522
rect 561971 312450 562017 312488
rect 561971 312416 561977 312450
rect 562011 312416 562017 312450
rect 561971 312378 562017 312416
rect 561971 312344 561977 312378
rect 562011 312344 562017 312378
rect 561971 312306 562017 312344
rect 561971 312272 561977 312306
rect 562011 312272 562017 312306
rect 561971 312234 562017 312272
rect 561971 312200 561977 312234
rect 562011 312200 562017 312234
rect 561971 312162 562017 312200
rect 561971 312128 561977 312162
rect 562011 312128 562017 312162
rect 561971 312090 562017 312128
rect 561971 312056 561977 312090
rect 562011 312056 562017 312090
rect 561971 312018 562017 312056
rect 561971 311984 561977 312018
rect 562011 311984 562017 312018
rect 561971 311946 562017 311984
rect 561971 311912 561977 311946
rect 562011 311912 562017 311946
rect 561971 311874 562017 311912
rect 561971 311840 561977 311874
rect 562011 311840 562017 311874
rect 561971 311802 562017 311840
rect 561971 311768 561977 311802
rect 562011 311768 562017 311802
rect 561971 311730 562017 311768
rect 561971 311696 561977 311730
rect 562011 311696 562017 311730
rect 561971 311681 562017 311696
rect 562229 312666 562275 312681
rect 562229 312632 562235 312666
rect 562269 312632 562275 312666
rect 562229 312594 562275 312632
rect 562229 312560 562235 312594
rect 562269 312560 562275 312594
rect 562229 312522 562275 312560
rect 562229 312488 562235 312522
rect 562269 312488 562275 312522
rect 562229 312450 562275 312488
rect 562229 312416 562235 312450
rect 562269 312416 562275 312450
rect 562229 312378 562275 312416
rect 562229 312344 562235 312378
rect 562269 312344 562275 312378
rect 562229 312306 562275 312344
rect 562229 312272 562235 312306
rect 562269 312272 562275 312306
rect 562229 312234 562275 312272
rect 562229 312200 562235 312234
rect 562269 312200 562275 312234
rect 562229 312162 562275 312200
rect 562229 312128 562235 312162
rect 562269 312128 562275 312162
rect 562229 312090 562275 312128
rect 562229 312056 562235 312090
rect 562269 312056 562275 312090
rect 562229 312018 562275 312056
rect 562229 311984 562235 312018
rect 562269 311984 562275 312018
rect 562229 311946 562275 311984
rect 562229 311912 562235 311946
rect 562269 311912 562275 311946
rect 562229 311874 562275 311912
rect 562229 311840 562235 311874
rect 562269 311840 562275 311874
rect 562229 311802 562275 311840
rect 562229 311768 562235 311802
rect 562269 311768 562275 311802
rect 562229 311730 562275 311768
rect 562229 311696 562235 311730
rect 562269 311696 562275 311730
rect 562229 311681 562275 311696
rect 562487 312666 562533 312681
rect 562487 312632 562493 312666
rect 562527 312632 562533 312666
rect 562487 312594 562533 312632
rect 562487 312560 562493 312594
rect 562527 312560 562533 312594
rect 562487 312522 562533 312560
rect 562487 312488 562493 312522
rect 562527 312488 562533 312522
rect 562487 312450 562533 312488
rect 562487 312416 562493 312450
rect 562527 312416 562533 312450
rect 562487 312378 562533 312416
rect 562487 312344 562493 312378
rect 562527 312344 562533 312378
rect 562487 312306 562533 312344
rect 562487 312272 562493 312306
rect 562527 312272 562533 312306
rect 562487 312234 562533 312272
rect 562487 312200 562493 312234
rect 562527 312200 562533 312234
rect 562487 312162 562533 312200
rect 562487 312128 562493 312162
rect 562527 312128 562533 312162
rect 562487 312090 562533 312128
rect 562487 312056 562493 312090
rect 562527 312056 562533 312090
rect 562487 312018 562533 312056
rect 562487 311984 562493 312018
rect 562527 311984 562533 312018
rect 562487 311946 562533 311984
rect 562487 311912 562493 311946
rect 562527 311912 562533 311946
rect 562487 311874 562533 311912
rect 562487 311840 562493 311874
rect 562527 311840 562533 311874
rect 562487 311802 562533 311840
rect 562487 311768 562493 311802
rect 562527 311768 562533 311802
rect 562487 311730 562533 311768
rect 562487 311696 562493 311730
rect 562527 311696 562533 311730
rect 562487 311681 562533 311696
rect 562745 312666 562791 312681
rect 562745 312632 562751 312666
rect 562785 312632 562791 312666
rect 562745 312594 562791 312632
rect 562745 312560 562751 312594
rect 562785 312560 562791 312594
rect 562745 312522 562791 312560
rect 562745 312488 562751 312522
rect 562785 312488 562791 312522
rect 562745 312450 562791 312488
rect 562745 312416 562751 312450
rect 562785 312416 562791 312450
rect 562745 312378 562791 312416
rect 562745 312344 562751 312378
rect 562785 312344 562791 312378
rect 562745 312306 562791 312344
rect 562745 312272 562751 312306
rect 562785 312272 562791 312306
rect 562745 312234 562791 312272
rect 562745 312200 562751 312234
rect 562785 312200 562791 312234
rect 562745 312162 562791 312200
rect 562745 312128 562751 312162
rect 562785 312128 562791 312162
rect 562745 312090 562791 312128
rect 562745 312056 562751 312090
rect 562785 312056 562791 312090
rect 562745 312018 562791 312056
rect 562745 311984 562751 312018
rect 562785 311984 562791 312018
rect 562745 311946 562791 311984
rect 562745 311912 562751 311946
rect 562785 311912 562791 311946
rect 562745 311874 562791 311912
rect 562745 311840 562751 311874
rect 562785 311840 562791 311874
rect 562745 311802 562791 311840
rect 562745 311768 562751 311802
rect 562785 311768 562791 311802
rect 562745 311730 562791 311768
rect 562745 311696 562751 311730
rect 562785 311696 562791 311730
rect 562745 311681 562791 311696
rect 563003 312666 563049 312681
rect 563003 312632 563009 312666
rect 563043 312632 563049 312666
rect 563003 312594 563049 312632
rect 563003 312560 563009 312594
rect 563043 312560 563049 312594
rect 563003 312522 563049 312560
rect 563003 312488 563009 312522
rect 563043 312488 563049 312522
rect 563003 312450 563049 312488
rect 563003 312416 563009 312450
rect 563043 312416 563049 312450
rect 563003 312378 563049 312416
rect 563003 312344 563009 312378
rect 563043 312344 563049 312378
rect 563003 312306 563049 312344
rect 563003 312272 563009 312306
rect 563043 312272 563049 312306
rect 563003 312234 563049 312272
rect 563003 312200 563009 312234
rect 563043 312200 563049 312234
rect 563003 312162 563049 312200
rect 563003 312128 563009 312162
rect 563043 312128 563049 312162
rect 563003 312090 563049 312128
rect 563003 312056 563009 312090
rect 563043 312056 563049 312090
rect 563003 312018 563049 312056
rect 563003 311984 563009 312018
rect 563043 311984 563049 312018
rect 563003 311946 563049 311984
rect 563003 311912 563009 311946
rect 563043 311912 563049 311946
rect 563003 311874 563049 311912
rect 563003 311840 563009 311874
rect 563043 311840 563049 311874
rect 563003 311802 563049 311840
rect 563003 311768 563009 311802
rect 563043 311768 563049 311802
rect 563003 311730 563049 311768
rect 563003 311696 563009 311730
rect 563043 311696 563049 311730
rect 563003 311681 563049 311696
rect 563261 312666 563307 312681
rect 563261 312632 563267 312666
rect 563301 312632 563307 312666
rect 563261 312594 563307 312632
rect 563261 312560 563267 312594
rect 563301 312560 563307 312594
rect 563261 312522 563307 312560
rect 563261 312488 563267 312522
rect 563301 312488 563307 312522
rect 563261 312450 563307 312488
rect 563261 312416 563267 312450
rect 563301 312416 563307 312450
rect 563261 312378 563307 312416
rect 563261 312344 563267 312378
rect 563301 312344 563307 312378
rect 563261 312306 563307 312344
rect 563261 312272 563267 312306
rect 563301 312272 563307 312306
rect 563261 312234 563307 312272
rect 563261 312200 563267 312234
rect 563301 312200 563307 312234
rect 563261 312162 563307 312200
rect 563261 312128 563267 312162
rect 563301 312128 563307 312162
rect 563261 312090 563307 312128
rect 563261 312056 563267 312090
rect 563301 312056 563307 312090
rect 563261 312018 563307 312056
rect 563261 311984 563267 312018
rect 563301 311984 563307 312018
rect 563261 311946 563307 311984
rect 563261 311912 563267 311946
rect 563301 311912 563307 311946
rect 563261 311874 563307 311912
rect 563261 311840 563267 311874
rect 563301 311840 563307 311874
rect 563261 311802 563307 311840
rect 563261 311768 563267 311802
rect 563301 311768 563307 311802
rect 563261 311730 563307 311768
rect 563261 311696 563267 311730
rect 563301 311696 563307 311730
rect 563261 311681 563307 311696
rect 563519 312666 563565 312681
rect 563519 312632 563525 312666
rect 563559 312632 563565 312666
rect 563519 312594 563565 312632
rect 563519 312560 563525 312594
rect 563559 312560 563565 312594
rect 563519 312522 563565 312560
rect 563519 312488 563525 312522
rect 563559 312488 563565 312522
rect 563519 312450 563565 312488
rect 563519 312416 563525 312450
rect 563559 312416 563565 312450
rect 563519 312378 563565 312416
rect 563519 312344 563525 312378
rect 563559 312344 563565 312378
rect 563519 312306 563565 312344
rect 563519 312272 563525 312306
rect 563559 312272 563565 312306
rect 563519 312234 563565 312272
rect 563519 312200 563525 312234
rect 563559 312200 563565 312234
rect 563519 312162 563565 312200
rect 563519 312128 563525 312162
rect 563559 312128 563565 312162
rect 563519 312090 563565 312128
rect 563519 312056 563525 312090
rect 563559 312056 563565 312090
rect 563519 312018 563565 312056
rect 563519 311984 563525 312018
rect 563559 311984 563565 312018
rect 563519 311946 563565 311984
rect 563519 311912 563525 311946
rect 563559 311912 563565 311946
rect 563519 311874 563565 311912
rect 563519 311840 563525 311874
rect 563559 311840 563565 311874
rect 563519 311802 563565 311840
rect 563519 311768 563525 311802
rect 563559 311768 563565 311802
rect 563519 311730 563565 311768
rect 563519 311696 563525 311730
rect 563559 311696 563565 311730
rect 563519 311681 563565 311696
rect 563777 312666 563823 312681
rect 563777 312632 563783 312666
rect 563817 312632 563823 312666
rect 563777 312594 563823 312632
rect 563777 312560 563783 312594
rect 563817 312560 563823 312594
rect 563777 312522 563823 312560
rect 563777 312488 563783 312522
rect 563817 312488 563823 312522
rect 563777 312450 563823 312488
rect 563777 312416 563783 312450
rect 563817 312416 563823 312450
rect 563777 312378 563823 312416
rect 563777 312344 563783 312378
rect 563817 312344 563823 312378
rect 563777 312306 563823 312344
rect 563777 312272 563783 312306
rect 563817 312272 563823 312306
rect 563777 312234 563823 312272
rect 563777 312200 563783 312234
rect 563817 312200 563823 312234
rect 563777 312162 563823 312200
rect 563777 312128 563783 312162
rect 563817 312128 563823 312162
rect 563777 312090 563823 312128
rect 563777 312056 563783 312090
rect 563817 312056 563823 312090
rect 563777 312018 563823 312056
rect 563777 311984 563783 312018
rect 563817 311984 563823 312018
rect 563777 311946 563823 311984
rect 563777 311912 563783 311946
rect 563817 311912 563823 311946
rect 563777 311874 563823 311912
rect 563777 311840 563783 311874
rect 563817 311840 563823 311874
rect 563777 311802 563823 311840
rect 563777 311768 563783 311802
rect 563817 311768 563823 311802
rect 563777 311730 563823 311768
rect 563777 311696 563783 311730
rect 563817 311696 563823 311730
rect 563777 311681 563823 311696
rect 564035 312666 564081 312681
rect 564035 312632 564041 312666
rect 564075 312632 564081 312666
rect 564035 312594 564081 312632
rect 564035 312560 564041 312594
rect 564075 312560 564081 312594
rect 564035 312522 564081 312560
rect 564035 312488 564041 312522
rect 564075 312488 564081 312522
rect 564035 312450 564081 312488
rect 564035 312416 564041 312450
rect 564075 312416 564081 312450
rect 564035 312378 564081 312416
rect 564035 312344 564041 312378
rect 564075 312344 564081 312378
rect 564035 312306 564081 312344
rect 564035 312272 564041 312306
rect 564075 312272 564081 312306
rect 564035 312234 564081 312272
rect 564035 312200 564041 312234
rect 564075 312200 564081 312234
rect 564035 312162 564081 312200
rect 564035 312128 564041 312162
rect 564075 312128 564081 312162
rect 564035 312090 564081 312128
rect 564035 312056 564041 312090
rect 564075 312056 564081 312090
rect 564035 312018 564081 312056
rect 564035 311984 564041 312018
rect 564075 311984 564081 312018
rect 564035 311946 564081 311984
rect 564035 311912 564041 311946
rect 564075 311912 564081 311946
rect 564035 311874 564081 311912
rect 564035 311840 564041 311874
rect 564075 311840 564081 311874
rect 564035 311802 564081 311840
rect 564035 311768 564041 311802
rect 564075 311768 564081 311802
rect 564035 311730 564081 311768
rect 564035 311696 564041 311730
rect 564075 311696 564081 311730
rect 564035 311681 564081 311696
rect 564293 312666 564339 312681
rect 564293 312632 564299 312666
rect 564333 312632 564339 312666
rect 564293 312594 564339 312632
rect 564293 312560 564299 312594
rect 564333 312560 564339 312594
rect 564293 312522 564339 312560
rect 564293 312488 564299 312522
rect 564333 312488 564339 312522
rect 564293 312450 564339 312488
rect 564293 312416 564299 312450
rect 564333 312416 564339 312450
rect 564293 312378 564339 312416
rect 564293 312344 564299 312378
rect 564333 312344 564339 312378
rect 564293 312306 564339 312344
rect 564293 312272 564299 312306
rect 564333 312272 564339 312306
rect 564293 312234 564339 312272
rect 564293 312200 564299 312234
rect 564333 312200 564339 312234
rect 564293 312162 564339 312200
rect 564293 312128 564299 312162
rect 564333 312128 564339 312162
rect 564293 312090 564339 312128
rect 564293 312056 564299 312090
rect 564333 312056 564339 312090
rect 564293 312018 564339 312056
rect 564293 311984 564299 312018
rect 564333 311984 564339 312018
rect 564293 311946 564339 311984
rect 564293 311912 564299 311946
rect 564333 311912 564339 311946
rect 564293 311874 564339 311912
rect 564293 311840 564299 311874
rect 564333 311840 564339 311874
rect 564293 311802 564339 311840
rect 564293 311768 564299 311802
rect 564333 311768 564339 311802
rect 564293 311730 564339 311768
rect 564293 311696 564299 311730
rect 564333 311696 564339 311730
rect 564293 311681 564339 311696
rect 564551 312666 564597 312681
rect 564551 312632 564557 312666
rect 564591 312632 564597 312666
rect 564551 312594 564597 312632
rect 564551 312560 564557 312594
rect 564591 312560 564597 312594
rect 564551 312522 564597 312560
rect 564551 312488 564557 312522
rect 564591 312488 564597 312522
rect 564551 312450 564597 312488
rect 564551 312416 564557 312450
rect 564591 312416 564597 312450
rect 564551 312378 564597 312416
rect 564551 312344 564557 312378
rect 564591 312344 564597 312378
rect 564551 312306 564597 312344
rect 564551 312272 564557 312306
rect 564591 312272 564597 312306
rect 564551 312234 564597 312272
rect 564551 312200 564557 312234
rect 564591 312200 564597 312234
rect 564551 312162 564597 312200
rect 564551 312128 564557 312162
rect 564591 312128 564597 312162
rect 564551 312090 564597 312128
rect 564551 312056 564557 312090
rect 564591 312056 564597 312090
rect 564551 312018 564597 312056
rect 564551 311984 564557 312018
rect 564591 311984 564597 312018
rect 564551 311946 564597 311984
rect 564551 311912 564557 311946
rect 564591 311912 564597 311946
rect 564551 311874 564597 311912
rect 564551 311840 564557 311874
rect 564591 311840 564597 311874
rect 564551 311802 564597 311840
rect 564551 311768 564557 311802
rect 564591 311768 564597 311802
rect 564551 311730 564597 311768
rect 564551 311696 564557 311730
rect 564591 311696 564597 311730
rect 564551 311681 564597 311696
rect 564809 312666 564855 312681
rect 564809 312632 564815 312666
rect 564849 312632 564855 312666
rect 564809 312594 564855 312632
rect 564809 312560 564815 312594
rect 564849 312560 564855 312594
rect 564809 312522 564855 312560
rect 564809 312488 564815 312522
rect 564849 312488 564855 312522
rect 564809 312450 564855 312488
rect 564809 312416 564815 312450
rect 564849 312416 564855 312450
rect 564809 312378 564855 312416
rect 564809 312344 564815 312378
rect 564849 312344 564855 312378
rect 564809 312306 564855 312344
rect 564809 312272 564815 312306
rect 564849 312272 564855 312306
rect 564809 312234 564855 312272
rect 564809 312200 564815 312234
rect 564849 312200 564855 312234
rect 564809 312162 564855 312200
rect 564809 312128 564815 312162
rect 564849 312128 564855 312162
rect 564809 312090 564855 312128
rect 564809 312056 564815 312090
rect 564849 312056 564855 312090
rect 564809 312018 564855 312056
rect 564809 311984 564815 312018
rect 564849 311984 564855 312018
rect 564809 311946 564855 311984
rect 564809 311912 564815 311946
rect 564849 311912 564855 311946
rect 564809 311874 564855 311912
rect 564809 311840 564815 311874
rect 564849 311840 564855 311874
rect 564809 311802 564855 311840
rect 564809 311768 564815 311802
rect 564849 311768 564855 311802
rect 564809 311730 564855 311768
rect 564809 311696 564815 311730
rect 564849 311696 564855 311730
rect 564809 311681 564855 311696
rect 565067 312666 565113 312681
rect 565067 312632 565073 312666
rect 565107 312632 565113 312666
rect 565067 312594 565113 312632
rect 565067 312560 565073 312594
rect 565107 312560 565113 312594
rect 565067 312522 565113 312560
rect 565067 312488 565073 312522
rect 565107 312488 565113 312522
rect 565067 312450 565113 312488
rect 565067 312416 565073 312450
rect 565107 312416 565113 312450
rect 565067 312378 565113 312416
rect 565067 312344 565073 312378
rect 565107 312344 565113 312378
rect 565067 312306 565113 312344
rect 565067 312272 565073 312306
rect 565107 312272 565113 312306
rect 565067 312234 565113 312272
rect 565067 312200 565073 312234
rect 565107 312200 565113 312234
rect 565067 312162 565113 312200
rect 565067 312128 565073 312162
rect 565107 312128 565113 312162
rect 565067 312090 565113 312128
rect 565067 312056 565073 312090
rect 565107 312056 565113 312090
rect 565067 312018 565113 312056
rect 565067 311984 565073 312018
rect 565107 311984 565113 312018
rect 565067 311946 565113 311984
rect 565067 311912 565073 311946
rect 565107 311912 565113 311946
rect 565067 311874 565113 311912
rect 565067 311840 565073 311874
rect 565107 311840 565113 311874
rect 565067 311802 565113 311840
rect 565067 311768 565073 311802
rect 565107 311768 565113 311802
rect 565067 311730 565113 311768
rect 565067 311696 565073 311730
rect 565107 311696 565113 311730
rect 565067 311681 565113 311696
rect 565325 312666 565371 312681
rect 565325 312632 565331 312666
rect 565365 312632 565371 312666
rect 565325 312594 565371 312632
rect 565325 312560 565331 312594
rect 565365 312560 565371 312594
rect 565325 312522 565371 312560
rect 565325 312488 565331 312522
rect 565365 312488 565371 312522
rect 565325 312450 565371 312488
rect 565325 312416 565331 312450
rect 565365 312416 565371 312450
rect 565325 312378 565371 312416
rect 565325 312344 565331 312378
rect 565365 312344 565371 312378
rect 565325 312306 565371 312344
rect 565325 312272 565331 312306
rect 565365 312272 565371 312306
rect 565325 312234 565371 312272
rect 565325 312200 565331 312234
rect 565365 312200 565371 312234
rect 565325 312162 565371 312200
rect 565325 312128 565331 312162
rect 565365 312128 565371 312162
rect 565325 312090 565371 312128
rect 565325 312056 565331 312090
rect 565365 312056 565371 312090
rect 565325 312018 565371 312056
rect 565325 311984 565331 312018
rect 565365 311984 565371 312018
rect 565325 311946 565371 311984
rect 565325 311912 565331 311946
rect 565365 311912 565371 311946
rect 565325 311874 565371 311912
rect 565325 311840 565331 311874
rect 565365 311840 565371 311874
rect 565325 311802 565371 311840
rect 565325 311768 565331 311802
rect 565365 311768 565371 311802
rect 565325 311730 565371 311768
rect 565325 311696 565331 311730
rect 565365 311696 565371 311730
rect 565325 311681 565371 311696
rect 565583 312666 565629 312681
rect 565583 312632 565589 312666
rect 565623 312632 565629 312666
rect 565583 312594 565629 312632
rect 565583 312560 565589 312594
rect 565623 312560 565629 312594
rect 565583 312522 565629 312560
rect 565583 312488 565589 312522
rect 565623 312488 565629 312522
rect 565583 312450 565629 312488
rect 565583 312416 565589 312450
rect 565623 312416 565629 312450
rect 565583 312378 565629 312416
rect 565583 312344 565589 312378
rect 565623 312344 565629 312378
rect 565583 312306 565629 312344
rect 565583 312272 565589 312306
rect 565623 312272 565629 312306
rect 565583 312234 565629 312272
rect 565583 312200 565589 312234
rect 565623 312200 565629 312234
rect 565583 312162 565629 312200
rect 565583 312128 565589 312162
rect 565623 312128 565629 312162
rect 565583 312090 565629 312128
rect 565583 312056 565589 312090
rect 565623 312056 565629 312090
rect 565583 312018 565629 312056
rect 565583 311984 565589 312018
rect 565623 311984 565629 312018
rect 565583 311946 565629 311984
rect 565583 311912 565589 311946
rect 565623 311912 565629 311946
rect 565583 311874 565629 311912
rect 565583 311840 565589 311874
rect 565623 311840 565629 311874
rect 565583 311802 565629 311840
rect 565583 311768 565589 311802
rect 565623 311768 565629 311802
rect 565583 311730 565629 311768
rect 565583 311696 565589 311730
rect 565623 311696 565629 311730
rect 565583 311681 565629 311696
rect 566130 311693 566376 313626
rect 573560 313191 573784 314307
rect 580858 313787 580962 313791
rect 580770 313779 580962 313787
rect 580762 313753 580968 313779
rect 580762 313637 580775 313753
rect 580955 313637 580968 313753
rect 580762 313611 580968 313637
rect 573560 313148 580492 313191
rect 573560 313114 575177 313148
rect 575211 313114 575377 313148
rect 575411 313114 575577 313148
rect 575611 313114 575777 313148
rect 575811 313114 575977 313148
rect 576011 313114 576177 313148
rect 576211 313114 576377 313148
rect 576411 313114 576577 313148
rect 576611 313114 576777 313148
rect 576811 313114 576977 313148
rect 577011 313114 577177 313148
rect 577211 313114 577377 313148
rect 577411 313114 577577 313148
rect 577611 313114 577777 313148
rect 577811 313114 577977 313148
rect 578011 313114 578177 313148
rect 578211 313114 578377 313148
rect 578411 313114 578577 313148
rect 578611 313114 578777 313148
rect 578811 313114 578977 313148
rect 579011 313114 579177 313148
rect 579211 313114 579377 313148
rect 579411 313114 579577 313148
rect 579611 313114 579777 313148
rect 579811 313114 579977 313148
rect 580011 313114 580177 313148
rect 580211 313114 580492 313148
rect 573560 313071 580492 313114
rect 573560 311751 573814 313071
rect 575147 312736 575193 312751
rect 575147 312702 575153 312736
rect 575187 312702 575193 312736
rect 575147 312664 575193 312702
rect 575147 312630 575153 312664
rect 575187 312630 575193 312664
rect 575147 312592 575193 312630
rect 575147 312558 575153 312592
rect 575187 312558 575193 312592
rect 575147 312520 575193 312558
rect 575147 312486 575153 312520
rect 575187 312486 575193 312520
rect 575147 312448 575193 312486
rect 575147 312414 575153 312448
rect 575187 312414 575193 312448
rect 575147 312376 575193 312414
rect 575147 312342 575153 312376
rect 575187 312342 575193 312376
rect 575147 312304 575193 312342
rect 575147 312270 575153 312304
rect 575187 312270 575193 312304
rect 575147 312232 575193 312270
rect 575147 312198 575153 312232
rect 575187 312198 575193 312232
rect 575147 312160 575193 312198
rect 575147 312126 575153 312160
rect 575187 312126 575193 312160
rect 575147 312088 575193 312126
rect 575147 312054 575153 312088
rect 575187 312054 575193 312088
rect 575147 312016 575193 312054
rect 575147 311982 575153 312016
rect 575187 311982 575193 312016
rect 575147 311944 575193 311982
rect 575147 311910 575153 311944
rect 575187 311910 575193 311944
rect 575147 311872 575193 311910
rect 575147 311838 575153 311872
rect 575187 311838 575193 311872
rect 575147 311800 575193 311838
rect 575147 311766 575153 311800
rect 575187 311766 575193 311800
rect 575147 311751 575193 311766
rect 575405 312736 575451 312751
rect 575405 312702 575411 312736
rect 575445 312702 575451 312736
rect 575405 312664 575451 312702
rect 575405 312630 575411 312664
rect 575445 312630 575451 312664
rect 575405 312592 575451 312630
rect 575405 312558 575411 312592
rect 575445 312558 575451 312592
rect 575405 312520 575451 312558
rect 575405 312486 575411 312520
rect 575445 312486 575451 312520
rect 575405 312448 575451 312486
rect 575405 312414 575411 312448
rect 575445 312414 575451 312448
rect 575405 312376 575451 312414
rect 575405 312342 575411 312376
rect 575445 312342 575451 312376
rect 575405 312304 575451 312342
rect 575405 312270 575411 312304
rect 575445 312270 575451 312304
rect 575405 312232 575451 312270
rect 575405 312198 575411 312232
rect 575445 312198 575451 312232
rect 575405 312160 575451 312198
rect 575405 312126 575411 312160
rect 575445 312126 575451 312160
rect 575405 312088 575451 312126
rect 575405 312054 575411 312088
rect 575445 312054 575451 312088
rect 575405 312016 575451 312054
rect 575405 311982 575411 312016
rect 575445 311982 575451 312016
rect 575405 311944 575451 311982
rect 575405 311910 575411 311944
rect 575445 311910 575451 311944
rect 575405 311872 575451 311910
rect 575405 311838 575411 311872
rect 575445 311838 575451 311872
rect 575405 311800 575451 311838
rect 575405 311766 575411 311800
rect 575445 311766 575451 311800
rect 575405 311751 575451 311766
rect 575663 312736 575709 312751
rect 575663 312702 575669 312736
rect 575703 312702 575709 312736
rect 575663 312664 575709 312702
rect 575663 312630 575669 312664
rect 575703 312630 575709 312664
rect 575663 312592 575709 312630
rect 575663 312558 575669 312592
rect 575703 312558 575709 312592
rect 575663 312520 575709 312558
rect 575663 312486 575669 312520
rect 575703 312486 575709 312520
rect 575663 312448 575709 312486
rect 575663 312414 575669 312448
rect 575703 312414 575709 312448
rect 575663 312376 575709 312414
rect 575663 312342 575669 312376
rect 575703 312342 575709 312376
rect 575663 312304 575709 312342
rect 575663 312270 575669 312304
rect 575703 312270 575709 312304
rect 575663 312232 575709 312270
rect 575663 312198 575669 312232
rect 575703 312198 575709 312232
rect 575663 312160 575709 312198
rect 575663 312126 575669 312160
rect 575703 312126 575709 312160
rect 575663 312088 575709 312126
rect 575663 312054 575669 312088
rect 575703 312054 575709 312088
rect 575663 312016 575709 312054
rect 575663 311982 575669 312016
rect 575703 311982 575709 312016
rect 575663 311944 575709 311982
rect 575663 311910 575669 311944
rect 575703 311910 575709 311944
rect 575663 311872 575709 311910
rect 575663 311838 575669 311872
rect 575703 311838 575709 311872
rect 575663 311800 575709 311838
rect 575663 311766 575669 311800
rect 575703 311766 575709 311800
rect 575663 311751 575709 311766
rect 575921 312736 575967 312751
rect 575921 312702 575927 312736
rect 575961 312702 575967 312736
rect 575921 312664 575967 312702
rect 575921 312630 575927 312664
rect 575961 312630 575967 312664
rect 575921 312592 575967 312630
rect 575921 312558 575927 312592
rect 575961 312558 575967 312592
rect 575921 312520 575967 312558
rect 575921 312486 575927 312520
rect 575961 312486 575967 312520
rect 575921 312448 575967 312486
rect 575921 312414 575927 312448
rect 575961 312414 575967 312448
rect 575921 312376 575967 312414
rect 575921 312342 575927 312376
rect 575961 312342 575967 312376
rect 575921 312304 575967 312342
rect 575921 312270 575927 312304
rect 575961 312270 575967 312304
rect 575921 312232 575967 312270
rect 575921 312198 575927 312232
rect 575961 312198 575967 312232
rect 575921 312160 575967 312198
rect 575921 312126 575927 312160
rect 575961 312126 575967 312160
rect 575921 312088 575967 312126
rect 575921 312054 575927 312088
rect 575961 312054 575967 312088
rect 575921 312016 575967 312054
rect 575921 311982 575927 312016
rect 575961 311982 575967 312016
rect 575921 311944 575967 311982
rect 575921 311910 575927 311944
rect 575961 311910 575967 311944
rect 575921 311872 575967 311910
rect 575921 311838 575927 311872
rect 575961 311838 575967 311872
rect 575921 311800 575967 311838
rect 575921 311766 575927 311800
rect 575961 311766 575967 311800
rect 575921 311751 575967 311766
rect 576179 312736 576225 312751
rect 576179 312702 576185 312736
rect 576219 312702 576225 312736
rect 576179 312664 576225 312702
rect 576179 312630 576185 312664
rect 576219 312630 576225 312664
rect 576179 312592 576225 312630
rect 576179 312558 576185 312592
rect 576219 312558 576225 312592
rect 576179 312520 576225 312558
rect 576179 312486 576185 312520
rect 576219 312486 576225 312520
rect 576179 312448 576225 312486
rect 576179 312414 576185 312448
rect 576219 312414 576225 312448
rect 576179 312376 576225 312414
rect 576179 312342 576185 312376
rect 576219 312342 576225 312376
rect 576179 312304 576225 312342
rect 576179 312270 576185 312304
rect 576219 312270 576225 312304
rect 576179 312232 576225 312270
rect 576179 312198 576185 312232
rect 576219 312198 576225 312232
rect 576179 312160 576225 312198
rect 576179 312126 576185 312160
rect 576219 312126 576225 312160
rect 576179 312088 576225 312126
rect 576179 312054 576185 312088
rect 576219 312054 576225 312088
rect 576179 312016 576225 312054
rect 576179 311982 576185 312016
rect 576219 311982 576225 312016
rect 576179 311944 576225 311982
rect 576179 311910 576185 311944
rect 576219 311910 576225 311944
rect 576179 311872 576225 311910
rect 576179 311838 576185 311872
rect 576219 311838 576225 311872
rect 576179 311800 576225 311838
rect 576179 311766 576185 311800
rect 576219 311766 576225 311800
rect 576179 311751 576225 311766
rect 576437 312736 576483 312751
rect 576437 312702 576443 312736
rect 576477 312702 576483 312736
rect 576437 312664 576483 312702
rect 576437 312630 576443 312664
rect 576477 312630 576483 312664
rect 576437 312592 576483 312630
rect 576437 312558 576443 312592
rect 576477 312558 576483 312592
rect 576437 312520 576483 312558
rect 576437 312486 576443 312520
rect 576477 312486 576483 312520
rect 576437 312448 576483 312486
rect 576437 312414 576443 312448
rect 576477 312414 576483 312448
rect 576437 312376 576483 312414
rect 576437 312342 576443 312376
rect 576477 312342 576483 312376
rect 576437 312304 576483 312342
rect 576437 312270 576443 312304
rect 576477 312270 576483 312304
rect 576437 312232 576483 312270
rect 576437 312198 576443 312232
rect 576477 312198 576483 312232
rect 576437 312160 576483 312198
rect 576437 312126 576443 312160
rect 576477 312126 576483 312160
rect 576437 312088 576483 312126
rect 576437 312054 576443 312088
rect 576477 312054 576483 312088
rect 576437 312016 576483 312054
rect 576437 311982 576443 312016
rect 576477 311982 576483 312016
rect 576437 311944 576483 311982
rect 576437 311910 576443 311944
rect 576477 311910 576483 311944
rect 576437 311872 576483 311910
rect 576437 311838 576443 311872
rect 576477 311838 576483 311872
rect 576437 311800 576483 311838
rect 576437 311766 576443 311800
rect 576477 311766 576483 311800
rect 576437 311751 576483 311766
rect 576695 312736 576741 312751
rect 576695 312702 576701 312736
rect 576735 312702 576741 312736
rect 576695 312664 576741 312702
rect 576695 312630 576701 312664
rect 576735 312630 576741 312664
rect 576695 312592 576741 312630
rect 576695 312558 576701 312592
rect 576735 312558 576741 312592
rect 576695 312520 576741 312558
rect 576695 312486 576701 312520
rect 576735 312486 576741 312520
rect 576695 312448 576741 312486
rect 576695 312414 576701 312448
rect 576735 312414 576741 312448
rect 576695 312376 576741 312414
rect 576695 312342 576701 312376
rect 576735 312342 576741 312376
rect 576695 312304 576741 312342
rect 576695 312270 576701 312304
rect 576735 312270 576741 312304
rect 576695 312232 576741 312270
rect 576695 312198 576701 312232
rect 576735 312198 576741 312232
rect 576695 312160 576741 312198
rect 576695 312126 576701 312160
rect 576735 312126 576741 312160
rect 576695 312088 576741 312126
rect 576695 312054 576701 312088
rect 576735 312054 576741 312088
rect 576695 312016 576741 312054
rect 576695 311982 576701 312016
rect 576735 311982 576741 312016
rect 576695 311944 576741 311982
rect 576695 311910 576701 311944
rect 576735 311910 576741 311944
rect 576695 311872 576741 311910
rect 576695 311838 576701 311872
rect 576735 311838 576741 311872
rect 576695 311800 576741 311838
rect 576695 311766 576701 311800
rect 576735 311766 576741 311800
rect 576695 311751 576741 311766
rect 576953 312736 576999 312751
rect 576953 312702 576959 312736
rect 576993 312702 576999 312736
rect 576953 312664 576999 312702
rect 576953 312630 576959 312664
rect 576993 312630 576999 312664
rect 576953 312592 576999 312630
rect 576953 312558 576959 312592
rect 576993 312558 576999 312592
rect 576953 312520 576999 312558
rect 576953 312486 576959 312520
rect 576993 312486 576999 312520
rect 576953 312448 576999 312486
rect 576953 312414 576959 312448
rect 576993 312414 576999 312448
rect 576953 312376 576999 312414
rect 576953 312342 576959 312376
rect 576993 312342 576999 312376
rect 576953 312304 576999 312342
rect 576953 312270 576959 312304
rect 576993 312270 576999 312304
rect 576953 312232 576999 312270
rect 576953 312198 576959 312232
rect 576993 312198 576999 312232
rect 576953 312160 576999 312198
rect 576953 312126 576959 312160
rect 576993 312126 576999 312160
rect 576953 312088 576999 312126
rect 576953 312054 576959 312088
rect 576993 312054 576999 312088
rect 576953 312016 576999 312054
rect 576953 311982 576959 312016
rect 576993 311982 576999 312016
rect 576953 311944 576999 311982
rect 576953 311910 576959 311944
rect 576993 311910 576999 311944
rect 576953 311872 576999 311910
rect 576953 311838 576959 311872
rect 576993 311838 576999 311872
rect 576953 311800 576999 311838
rect 576953 311766 576959 311800
rect 576993 311766 576999 311800
rect 576953 311751 576999 311766
rect 577211 312736 577257 312751
rect 577211 312702 577217 312736
rect 577251 312702 577257 312736
rect 577211 312664 577257 312702
rect 577211 312630 577217 312664
rect 577251 312630 577257 312664
rect 577211 312592 577257 312630
rect 577211 312558 577217 312592
rect 577251 312558 577257 312592
rect 577211 312520 577257 312558
rect 577211 312486 577217 312520
rect 577251 312486 577257 312520
rect 577211 312448 577257 312486
rect 577211 312414 577217 312448
rect 577251 312414 577257 312448
rect 577211 312376 577257 312414
rect 577211 312342 577217 312376
rect 577251 312342 577257 312376
rect 577211 312304 577257 312342
rect 577211 312270 577217 312304
rect 577251 312270 577257 312304
rect 577211 312232 577257 312270
rect 577211 312198 577217 312232
rect 577251 312198 577257 312232
rect 577211 312160 577257 312198
rect 577211 312126 577217 312160
rect 577251 312126 577257 312160
rect 577211 312088 577257 312126
rect 577211 312054 577217 312088
rect 577251 312054 577257 312088
rect 577211 312016 577257 312054
rect 577211 311982 577217 312016
rect 577251 311982 577257 312016
rect 577211 311944 577257 311982
rect 577211 311910 577217 311944
rect 577251 311910 577257 311944
rect 577211 311872 577257 311910
rect 577211 311838 577217 311872
rect 577251 311838 577257 311872
rect 577211 311800 577257 311838
rect 577211 311766 577217 311800
rect 577251 311766 577257 311800
rect 577211 311751 577257 311766
rect 577469 312736 577515 312751
rect 577469 312702 577475 312736
rect 577509 312702 577515 312736
rect 577469 312664 577515 312702
rect 577469 312630 577475 312664
rect 577509 312630 577515 312664
rect 577469 312592 577515 312630
rect 577469 312558 577475 312592
rect 577509 312558 577515 312592
rect 577469 312520 577515 312558
rect 577469 312486 577475 312520
rect 577509 312486 577515 312520
rect 577469 312448 577515 312486
rect 577469 312414 577475 312448
rect 577509 312414 577515 312448
rect 577469 312376 577515 312414
rect 577469 312342 577475 312376
rect 577509 312342 577515 312376
rect 577469 312304 577515 312342
rect 577469 312270 577475 312304
rect 577509 312270 577515 312304
rect 577469 312232 577515 312270
rect 577469 312198 577475 312232
rect 577509 312198 577515 312232
rect 577469 312160 577515 312198
rect 577469 312126 577475 312160
rect 577509 312126 577515 312160
rect 577469 312088 577515 312126
rect 577469 312054 577475 312088
rect 577509 312054 577515 312088
rect 577469 312016 577515 312054
rect 577469 311982 577475 312016
rect 577509 311982 577515 312016
rect 577469 311944 577515 311982
rect 577469 311910 577475 311944
rect 577509 311910 577515 311944
rect 577469 311872 577515 311910
rect 577469 311838 577475 311872
rect 577509 311838 577515 311872
rect 577469 311800 577515 311838
rect 577469 311766 577475 311800
rect 577509 311766 577515 311800
rect 577469 311751 577515 311766
rect 577727 312736 577773 312751
rect 577727 312702 577733 312736
rect 577767 312702 577773 312736
rect 577727 312664 577773 312702
rect 577727 312630 577733 312664
rect 577767 312630 577773 312664
rect 577727 312592 577773 312630
rect 577727 312558 577733 312592
rect 577767 312558 577773 312592
rect 577727 312520 577773 312558
rect 577727 312486 577733 312520
rect 577767 312486 577773 312520
rect 577727 312448 577773 312486
rect 577727 312414 577733 312448
rect 577767 312414 577773 312448
rect 577727 312376 577773 312414
rect 577727 312342 577733 312376
rect 577767 312342 577773 312376
rect 577727 312304 577773 312342
rect 577727 312270 577733 312304
rect 577767 312270 577773 312304
rect 577727 312232 577773 312270
rect 577727 312198 577733 312232
rect 577767 312198 577773 312232
rect 577727 312160 577773 312198
rect 577727 312126 577733 312160
rect 577767 312126 577773 312160
rect 577727 312088 577773 312126
rect 577727 312054 577733 312088
rect 577767 312054 577773 312088
rect 577727 312016 577773 312054
rect 577727 311982 577733 312016
rect 577767 311982 577773 312016
rect 577727 311944 577773 311982
rect 577727 311910 577733 311944
rect 577767 311910 577773 311944
rect 577727 311872 577773 311910
rect 577727 311838 577733 311872
rect 577767 311838 577773 311872
rect 577727 311800 577773 311838
rect 577727 311766 577733 311800
rect 577767 311766 577773 311800
rect 577727 311751 577773 311766
rect 577985 312736 578031 312751
rect 577985 312702 577991 312736
rect 578025 312702 578031 312736
rect 577985 312664 578031 312702
rect 577985 312630 577991 312664
rect 578025 312630 578031 312664
rect 577985 312592 578031 312630
rect 577985 312558 577991 312592
rect 578025 312558 578031 312592
rect 577985 312520 578031 312558
rect 577985 312486 577991 312520
rect 578025 312486 578031 312520
rect 577985 312448 578031 312486
rect 577985 312414 577991 312448
rect 578025 312414 578031 312448
rect 577985 312376 578031 312414
rect 577985 312342 577991 312376
rect 578025 312342 578031 312376
rect 577985 312304 578031 312342
rect 577985 312270 577991 312304
rect 578025 312270 578031 312304
rect 577985 312232 578031 312270
rect 577985 312198 577991 312232
rect 578025 312198 578031 312232
rect 577985 312160 578031 312198
rect 577985 312126 577991 312160
rect 578025 312126 578031 312160
rect 577985 312088 578031 312126
rect 577985 312054 577991 312088
rect 578025 312054 578031 312088
rect 577985 312016 578031 312054
rect 577985 311982 577991 312016
rect 578025 311982 578031 312016
rect 577985 311944 578031 311982
rect 577985 311910 577991 311944
rect 578025 311910 578031 311944
rect 577985 311872 578031 311910
rect 577985 311838 577991 311872
rect 578025 311838 578031 311872
rect 577985 311800 578031 311838
rect 577985 311766 577991 311800
rect 578025 311766 578031 311800
rect 577985 311751 578031 311766
rect 578243 312736 578289 312751
rect 578243 312702 578249 312736
rect 578283 312702 578289 312736
rect 578243 312664 578289 312702
rect 578243 312630 578249 312664
rect 578283 312630 578289 312664
rect 578243 312592 578289 312630
rect 578243 312558 578249 312592
rect 578283 312558 578289 312592
rect 578243 312520 578289 312558
rect 578243 312486 578249 312520
rect 578283 312486 578289 312520
rect 578243 312448 578289 312486
rect 578243 312414 578249 312448
rect 578283 312414 578289 312448
rect 578243 312376 578289 312414
rect 578243 312342 578249 312376
rect 578283 312342 578289 312376
rect 578243 312304 578289 312342
rect 578243 312270 578249 312304
rect 578283 312270 578289 312304
rect 578243 312232 578289 312270
rect 578243 312198 578249 312232
rect 578283 312198 578289 312232
rect 578243 312160 578289 312198
rect 578243 312126 578249 312160
rect 578283 312126 578289 312160
rect 578243 312088 578289 312126
rect 578243 312054 578249 312088
rect 578283 312054 578289 312088
rect 578243 312016 578289 312054
rect 578243 311982 578249 312016
rect 578283 311982 578289 312016
rect 578243 311944 578289 311982
rect 578243 311910 578249 311944
rect 578283 311910 578289 311944
rect 578243 311872 578289 311910
rect 578243 311838 578249 311872
rect 578283 311838 578289 311872
rect 578243 311800 578289 311838
rect 578243 311766 578249 311800
rect 578283 311766 578289 311800
rect 578243 311751 578289 311766
rect 578501 312736 578547 312751
rect 578501 312702 578507 312736
rect 578541 312702 578547 312736
rect 578501 312664 578547 312702
rect 578501 312630 578507 312664
rect 578541 312630 578547 312664
rect 578501 312592 578547 312630
rect 578501 312558 578507 312592
rect 578541 312558 578547 312592
rect 578501 312520 578547 312558
rect 578501 312486 578507 312520
rect 578541 312486 578547 312520
rect 578501 312448 578547 312486
rect 578501 312414 578507 312448
rect 578541 312414 578547 312448
rect 578501 312376 578547 312414
rect 578501 312342 578507 312376
rect 578541 312342 578547 312376
rect 578501 312304 578547 312342
rect 578501 312270 578507 312304
rect 578541 312270 578547 312304
rect 578501 312232 578547 312270
rect 578501 312198 578507 312232
rect 578541 312198 578547 312232
rect 578501 312160 578547 312198
rect 578501 312126 578507 312160
rect 578541 312126 578547 312160
rect 578501 312088 578547 312126
rect 578501 312054 578507 312088
rect 578541 312054 578547 312088
rect 578501 312016 578547 312054
rect 578501 311982 578507 312016
rect 578541 311982 578547 312016
rect 578501 311944 578547 311982
rect 578501 311910 578507 311944
rect 578541 311910 578547 311944
rect 578501 311872 578547 311910
rect 578501 311838 578507 311872
rect 578541 311838 578547 311872
rect 578501 311800 578547 311838
rect 578501 311766 578507 311800
rect 578541 311766 578547 311800
rect 578501 311751 578547 311766
rect 578759 312736 578805 312751
rect 578759 312702 578765 312736
rect 578799 312702 578805 312736
rect 578759 312664 578805 312702
rect 578759 312630 578765 312664
rect 578799 312630 578805 312664
rect 578759 312592 578805 312630
rect 578759 312558 578765 312592
rect 578799 312558 578805 312592
rect 578759 312520 578805 312558
rect 578759 312486 578765 312520
rect 578799 312486 578805 312520
rect 578759 312448 578805 312486
rect 578759 312414 578765 312448
rect 578799 312414 578805 312448
rect 578759 312376 578805 312414
rect 578759 312342 578765 312376
rect 578799 312342 578805 312376
rect 578759 312304 578805 312342
rect 578759 312270 578765 312304
rect 578799 312270 578805 312304
rect 578759 312232 578805 312270
rect 578759 312198 578765 312232
rect 578799 312198 578805 312232
rect 578759 312160 578805 312198
rect 578759 312126 578765 312160
rect 578799 312126 578805 312160
rect 578759 312088 578805 312126
rect 578759 312054 578765 312088
rect 578799 312054 578805 312088
rect 578759 312016 578805 312054
rect 578759 311982 578765 312016
rect 578799 311982 578805 312016
rect 578759 311944 578805 311982
rect 578759 311910 578765 311944
rect 578799 311910 578805 311944
rect 578759 311872 578805 311910
rect 578759 311838 578765 311872
rect 578799 311838 578805 311872
rect 578759 311800 578805 311838
rect 578759 311766 578765 311800
rect 578799 311766 578805 311800
rect 578759 311751 578805 311766
rect 579017 312736 579063 312751
rect 579017 312702 579023 312736
rect 579057 312702 579063 312736
rect 579017 312664 579063 312702
rect 579017 312630 579023 312664
rect 579057 312630 579063 312664
rect 579017 312592 579063 312630
rect 579017 312558 579023 312592
rect 579057 312558 579063 312592
rect 579017 312520 579063 312558
rect 579017 312486 579023 312520
rect 579057 312486 579063 312520
rect 579017 312448 579063 312486
rect 579017 312414 579023 312448
rect 579057 312414 579063 312448
rect 579017 312376 579063 312414
rect 579017 312342 579023 312376
rect 579057 312342 579063 312376
rect 579017 312304 579063 312342
rect 579017 312270 579023 312304
rect 579057 312270 579063 312304
rect 579017 312232 579063 312270
rect 579017 312198 579023 312232
rect 579057 312198 579063 312232
rect 579017 312160 579063 312198
rect 579017 312126 579023 312160
rect 579057 312126 579063 312160
rect 579017 312088 579063 312126
rect 579017 312054 579023 312088
rect 579057 312054 579063 312088
rect 579017 312016 579063 312054
rect 579017 311982 579023 312016
rect 579057 311982 579063 312016
rect 579017 311944 579063 311982
rect 579017 311910 579023 311944
rect 579057 311910 579063 311944
rect 579017 311872 579063 311910
rect 579017 311838 579023 311872
rect 579057 311838 579063 311872
rect 579017 311800 579063 311838
rect 579017 311766 579023 311800
rect 579057 311766 579063 311800
rect 579017 311751 579063 311766
rect 579275 312736 579321 312751
rect 579275 312702 579281 312736
rect 579315 312702 579321 312736
rect 579275 312664 579321 312702
rect 579275 312630 579281 312664
rect 579315 312630 579321 312664
rect 579275 312592 579321 312630
rect 579275 312558 579281 312592
rect 579315 312558 579321 312592
rect 579275 312520 579321 312558
rect 579275 312486 579281 312520
rect 579315 312486 579321 312520
rect 579275 312448 579321 312486
rect 579275 312414 579281 312448
rect 579315 312414 579321 312448
rect 579275 312376 579321 312414
rect 579275 312342 579281 312376
rect 579315 312342 579321 312376
rect 579275 312304 579321 312342
rect 579275 312270 579281 312304
rect 579315 312270 579321 312304
rect 579275 312232 579321 312270
rect 579275 312198 579281 312232
rect 579315 312198 579321 312232
rect 579275 312160 579321 312198
rect 579275 312126 579281 312160
rect 579315 312126 579321 312160
rect 579275 312088 579321 312126
rect 579275 312054 579281 312088
rect 579315 312054 579321 312088
rect 579275 312016 579321 312054
rect 579275 311982 579281 312016
rect 579315 311982 579321 312016
rect 579275 311944 579321 311982
rect 579275 311910 579281 311944
rect 579315 311910 579321 311944
rect 579275 311872 579321 311910
rect 579275 311838 579281 311872
rect 579315 311838 579321 311872
rect 579275 311800 579321 311838
rect 579275 311766 579281 311800
rect 579315 311766 579321 311800
rect 579275 311751 579321 311766
rect 579533 312736 579579 312751
rect 579533 312702 579539 312736
rect 579573 312702 579579 312736
rect 579533 312664 579579 312702
rect 579533 312630 579539 312664
rect 579573 312630 579579 312664
rect 579533 312592 579579 312630
rect 579533 312558 579539 312592
rect 579573 312558 579579 312592
rect 579533 312520 579579 312558
rect 579533 312486 579539 312520
rect 579573 312486 579579 312520
rect 579533 312448 579579 312486
rect 579533 312414 579539 312448
rect 579573 312414 579579 312448
rect 579533 312376 579579 312414
rect 579533 312342 579539 312376
rect 579573 312342 579579 312376
rect 579533 312304 579579 312342
rect 579533 312270 579539 312304
rect 579573 312270 579579 312304
rect 579533 312232 579579 312270
rect 579533 312198 579539 312232
rect 579573 312198 579579 312232
rect 579533 312160 579579 312198
rect 579533 312126 579539 312160
rect 579573 312126 579579 312160
rect 579533 312088 579579 312126
rect 579533 312054 579539 312088
rect 579573 312054 579579 312088
rect 579533 312016 579579 312054
rect 579533 311982 579539 312016
rect 579573 311982 579579 312016
rect 579533 311944 579579 311982
rect 579533 311910 579539 311944
rect 579573 311910 579579 311944
rect 579533 311872 579579 311910
rect 579533 311838 579539 311872
rect 579573 311838 579579 311872
rect 579533 311800 579579 311838
rect 579533 311766 579539 311800
rect 579573 311766 579579 311800
rect 579533 311751 579579 311766
rect 579791 312736 579837 312751
rect 579791 312702 579797 312736
rect 579831 312702 579837 312736
rect 579791 312664 579837 312702
rect 579791 312630 579797 312664
rect 579831 312630 579837 312664
rect 579791 312592 579837 312630
rect 579791 312558 579797 312592
rect 579831 312558 579837 312592
rect 579791 312520 579837 312558
rect 579791 312486 579797 312520
rect 579831 312486 579837 312520
rect 579791 312448 579837 312486
rect 579791 312414 579797 312448
rect 579831 312414 579837 312448
rect 579791 312376 579837 312414
rect 579791 312342 579797 312376
rect 579831 312342 579837 312376
rect 579791 312304 579837 312342
rect 579791 312270 579797 312304
rect 579831 312270 579837 312304
rect 579791 312232 579837 312270
rect 579791 312198 579797 312232
rect 579831 312198 579837 312232
rect 579791 312160 579837 312198
rect 579791 312126 579797 312160
rect 579831 312126 579837 312160
rect 579791 312088 579837 312126
rect 579791 312054 579797 312088
rect 579831 312054 579837 312088
rect 579791 312016 579837 312054
rect 579791 311982 579797 312016
rect 579831 311982 579837 312016
rect 579791 311944 579837 311982
rect 579791 311910 579797 311944
rect 579831 311910 579837 311944
rect 579791 311872 579837 311910
rect 579791 311838 579797 311872
rect 579831 311838 579837 311872
rect 579791 311800 579837 311838
rect 579791 311766 579797 311800
rect 579831 311766 579837 311800
rect 579791 311751 579837 311766
rect 580049 312736 580095 312751
rect 580049 312702 580055 312736
rect 580089 312702 580095 312736
rect 580049 312664 580095 312702
rect 580049 312630 580055 312664
rect 580089 312630 580095 312664
rect 580049 312592 580095 312630
rect 580049 312558 580055 312592
rect 580089 312558 580095 312592
rect 580049 312520 580095 312558
rect 580049 312486 580055 312520
rect 580089 312486 580095 312520
rect 580049 312448 580095 312486
rect 580049 312414 580055 312448
rect 580089 312414 580095 312448
rect 580049 312376 580095 312414
rect 580049 312342 580055 312376
rect 580089 312342 580095 312376
rect 580049 312304 580095 312342
rect 580049 312270 580055 312304
rect 580089 312270 580095 312304
rect 580049 312232 580095 312270
rect 580049 312198 580055 312232
rect 580089 312198 580095 312232
rect 580049 312160 580095 312198
rect 580049 312126 580055 312160
rect 580089 312126 580095 312160
rect 580049 312088 580095 312126
rect 580049 312054 580055 312088
rect 580089 312054 580095 312088
rect 580049 312016 580095 312054
rect 580049 311982 580055 312016
rect 580089 311982 580095 312016
rect 580049 311944 580095 311982
rect 580049 311910 580055 311944
rect 580089 311910 580095 311944
rect 580049 311872 580095 311910
rect 580049 311838 580055 311872
rect 580089 311838 580095 311872
rect 580049 311800 580095 311838
rect 580049 311766 580055 311800
rect 580089 311766 580095 311800
rect 580049 311751 580095 311766
rect 580307 312736 580353 312751
rect 580307 312702 580313 312736
rect 580347 312702 580353 312736
rect 580307 312664 580353 312702
rect 580307 312630 580313 312664
rect 580347 312630 580353 312664
rect 580307 312592 580353 312630
rect 580307 312558 580313 312592
rect 580347 312558 580353 312592
rect 580307 312520 580353 312558
rect 580307 312486 580313 312520
rect 580347 312486 580353 312520
rect 580307 312448 580353 312486
rect 580307 312414 580313 312448
rect 580347 312414 580353 312448
rect 580307 312376 580353 312414
rect 580307 312342 580313 312376
rect 580347 312342 580353 312376
rect 580307 312304 580353 312342
rect 580307 312270 580313 312304
rect 580347 312270 580353 312304
rect 580307 312232 580353 312270
rect 580307 312198 580313 312232
rect 580347 312198 580353 312232
rect 580307 312160 580353 312198
rect 580307 312126 580313 312160
rect 580347 312126 580353 312160
rect 580307 312088 580353 312126
rect 580307 312054 580313 312088
rect 580347 312054 580353 312088
rect 580307 312016 580353 312054
rect 580307 311982 580313 312016
rect 580347 311982 580353 312016
rect 580307 311944 580353 311982
rect 580307 311910 580313 311944
rect 580347 311910 580353 311944
rect 580307 311872 580353 311910
rect 580307 311838 580313 311872
rect 580347 311838 580353 311872
rect 580307 311800 580353 311838
rect 580307 311766 580313 311800
rect 580347 311766 580353 311800
rect 580307 311751 580353 311766
rect 559860 311559 560254 311595
rect 559656 311545 560254 311559
rect 565826 311668 566376 311693
rect 565826 311562 565869 311668
rect 565975 311562 566376 311668
rect 565826 311545 566376 311562
rect 573446 311691 574060 311751
rect 559662 311241 559894 311545
rect 573446 311447 573523 311691
rect 573831 311599 574060 311691
rect 580770 311667 580962 313611
rect 580466 311628 580962 311667
rect 573831 311533 574966 311599
rect 580466 311594 580506 311628
rect 580540 311594 580962 311628
rect 580466 311563 580962 311594
rect 580466 311561 580580 311563
rect 573831 311486 574970 311533
rect 573831 311452 574899 311486
rect 574933 311452 574970 311486
rect 573831 311447 574970 311452
rect 573446 311405 574970 311447
rect 573446 311401 574966 311405
rect 573446 311391 574064 311401
rect 575106 311268 580492 311311
rect 559662 311198 565732 311241
rect 559662 311164 560617 311198
rect 560651 311164 560817 311198
rect 560851 311164 561017 311198
rect 561051 311164 561217 311198
rect 561251 311164 561417 311198
rect 561451 311164 561617 311198
rect 561651 311164 561817 311198
rect 561851 311164 562017 311198
rect 562051 311164 562217 311198
rect 562251 311164 562417 311198
rect 562451 311164 562617 311198
rect 562651 311164 562817 311198
rect 562851 311164 563017 311198
rect 563051 311164 563217 311198
rect 563251 311164 563417 311198
rect 563451 311164 563617 311198
rect 563651 311164 563817 311198
rect 563851 311164 564017 311198
rect 564051 311164 564217 311198
rect 564251 311164 564417 311198
rect 564451 311164 564617 311198
rect 564651 311164 564817 311198
rect 564851 311164 565017 311198
rect 565051 311164 565217 311198
rect 565251 311164 565417 311198
rect 565451 311181 565732 311198
rect 575106 311234 575177 311268
rect 575211 311234 575377 311268
rect 575411 311234 575577 311268
rect 575611 311234 575777 311268
rect 575811 311234 575977 311268
rect 576011 311234 576177 311268
rect 576211 311234 576377 311268
rect 576411 311234 576577 311268
rect 576611 311234 576777 311268
rect 576811 311234 576977 311268
rect 577011 311234 577177 311268
rect 577211 311234 577377 311268
rect 577411 311234 577577 311268
rect 577611 311234 577777 311268
rect 577811 311234 577977 311268
rect 578011 311234 578177 311268
rect 578211 311234 578377 311268
rect 578411 311234 578577 311268
rect 578611 311234 578777 311268
rect 578811 311234 578977 311268
rect 579011 311234 579177 311268
rect 579211 311234 579377 311268
rect 579411 311234 579577 311268
rect 579611 311234 579777 311268
rect 579811 311234 579977 311268
rect 580011 311234 580177 311268
rect 580211 311234 580492 311268
rect 575106 311191 580492 311234
rect 575106 311181 575364 311191
rect 565451 311164 575364 311181
rect 559662 311061 575364 311164
<< via1 >>
rect 566221 494137 566401 494317
rect 559831 492349 560011 492529
rect 580872 494161 581052 494341
rect 573579 491911 573887 492155
rect 566283 405286 566463 405466
rect 559755 403231 559935 403347
rect 580116 405330 580168 405382
rect 573462 402962 573824 403244
rect 566311 359801 566491 359981
rect 559740 357867 559920 358047
rect 580293 359861 580345 359913
rect 580293 359797 580345 359849
rect 573569 357612 573877 357920
rect 508620 356429 508736 356609
rect 566160 313626 566340 313806
rect 559680 311559 559860 311739
rect 580775 313637 580955 313753
rect 573523 311447 573831 311691
<< metal2 >>
rect 580870 494341 581054 494367
rect 566200 494317 566422 494329
rect 566200 494295 566221 494317
rect 566401 494295 566422 494317
rect 566200 494159 566203 494295
rect 566419 494159 566422 494295
rect 566200 494137 566221 494159
rect 566401 494137 566422 494159
rect 566200 494125 566422 494137
rect 580870 494161 580872 494341
rect 581052 494161 581054 494341
rect 580870 494135 581054 494161
rect 559816 492529 560026 492555
rect 559816 492349 559831 492529
rect 560011 492349 560026 492529
rect 559816 492323 560026 492349
rect 573578 492155 573888 492179
rect 573578 491911 573579 492155
rect 573887 491911 573888 492155
rect 573578 491887 573888 491911
rect 566270 405484 566476 405495
rect 566270 405466 566305 405484
rect 566441 405466 566476 405484
rect 566270 405286 566283 405466
rect 566463 405286 566476 405466
rect 580088 405384 580196 405421
rect 580088 405328 580114 405384
rect 580170 405328 580196 405384
rect 580088 405291 580196 405328
rect 566270 405268 566305 405286
rect 566441 405268 566476 405286
rect 566270 405257 566476 405268
rect 559750 403357 559940 403387
rect 559750 403347 559777 403357
rect 559913 403347 559940 403357
rect 559750 403231 559755 403347
rect 559935 403231 559940 403347
rect 559750 403221 559777 403231
rect 559913 403221 559940 403231
rect 559750 403191 559940 403221
rect 573462 403244 573824 403254
rect 573462 402952 573824 402962
rect 541978 389509 542092 389529
rect 541978 389453 542007 389509
rect 542063 389453 542092 389509
rect 541978 389433 542092 389453
rect 541972 380673 542094 380687
rect 541972 380617 542005 380673
rect 542061 380617 542094 380673
rect 541972 380593 542094 380617
rect 541972 380537 542005 380593
rect 542061 380537 542094 380593
rect 541972 380523 542094 380537
rect 566288 359981 566514 359997
rect 566288 359959 566311 359981
rect 566491 359959 566514 359981
rect 566288 359823 566293 359959
rect 566509 359823 566514 359959
rect 566288 359801 566311 359823
rect 566491 359801 566514 359823
rect 566288 359785 566514 359801
rect 580266 359913 580372 359925
rect 580266 359883 580293 359913
rect 580345 359883 580372 359913
rect 580266 359827 580291 359883
rect 580347 359827 580372 359883
rect 580266 359797 580293 359827
rect 580345 359797 580372 359827
rect 580266 359785 580372 359797
rect 559726 358047 559934 358071
rect 559726 357867 559740 358047
rect 559920 357867 559934 358047
rect 559726 357843 559934 357867
rect 573554 357920 573892 357939
rect 573554 357612 573569 357920
rect 573877 357612 573892 357920
rect 573554 357593 573892 357612
rect 508610 356609 508746 356621
rect 508610 356587 508620 356609
rect 508736 356587 508746 356609
rect 508610 356429 508620 356451
rect 508736 356429 508746 356451
rect 508610 356417 508746 356429
rect 566140 313806 566360 313823
rect 566140 313784 566160 313806
rect 566340 313784 566360 313806
rect 566140 313648 566142 313784
rect 566358 313648 566360 313784
rect 566140 313626 566160 313648
rect 566340 313626 566360 313648
rect 566140 313609 566360 313626
rect 580772 313763 580958 313789
rect 580772 313753 580797 313763
rect 580933 313753 580958 313763
rect 580772 313637 580775 313753
rect 580955 313637 580958 313753
rect 580772 313627 580797 313637
rect 580933 313627 580958 313637
rect 580772 313601 580958 313627
rect 559666 311739 559874 311763
rect 559666 311559 559680 311739
rect 559860 311559 559874 311739
rect 559666 311535 559874 311559
rect 573506 311691 573848 311719
rect 573506 311447 573523 311691
rect 573831 311447 573848 311691
rect 573506 311419 573848 311447
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 566203 494159 566221 494295
rect 566221 494159 566401 494295
rect 566401 494159 566419 494295
rect 580894 494183 581030 494319
rect 559853 492371 559989 492507
rect 573585 491925 573881 492141
rect 566305 405466 566441 405484
rect 566305 405286 566441 405466
rect 580114 405382 580170 405384
rect 580114 405330 580116 405382
rect 580116 405330 580168 405382
rect 580168 405330 580170 405382
rect 580114 405328 580170 405330
rect 566305 405268 566441 405286
rect 559777 403347 559913 403357
rect 559777 403231 559913 403347
rect 559777 403221 559913 403231
rect 573462 402962 573824 403244
rect 542007 389453 542063 389509
rect 542005 380617 542061 380673
rect 542005 380537 542061 380593
rect 566293 359823 566311 359959
rect 566311 359823 566491 359959
rect 566491 359823 566509 359959
rect 580291 359861 580293 359883
rect 580293 359861 580345 359883
rect 580345 359861 580347 359883
rect 580291 359849 580347 359861
rect 580291 359827 580293 359849
rect 580293 359827 580345 359849
rect 580345 359827 580347 359849
rect 559762 357889 559898 358025
rect 573575 357618 573871 357914
rect 508610 356451 508620 356587
rect 508620 356451 508736 356587
rect 508736 356451 508746 356587
rect 566142 313648 566160 313784
rect 566160 313648 566340 313784
rect 566340 313648 566358 313784
rect 580797 313753 580933 313763
rect 580797 313637 580933 313753
rect 580797 313627 580933 313637
rect 559702 311581 559838 311717
rect 573529 311461 573825 311677
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 703613 515394 704800
rect 510574 701285 515408 703613
rect 520594 703131 525394 704800
rect 510566 701189 515408 701285
rect 510566 700101 515400 701189
rect 510566 699273 515406 700101
rect 510552 697677 515406 699273
rect 510552 697351 515386 697677
rect 510552 696849 510735 697351
rect 510574 689927 510735 696849
rect 515199 689927 515386 697351
rect 510574 689675 515386 689927
rect 520568 697327 525402 703131
rect 566594 702300 571594 704800
rect 520568 689903 520735 697327
rect 525199 689903 525402 697327
rect 520568 689736 525402 689903
rect -800 680242 1700 685242
rect 582300 677984 584800 682984
rect -800 643842 1660 648642
rect 567119 644605 581246 644615
rect 567119 644584 582932 644605
rect 567119 644323 584800 644584
rect 567119 640099 567336 644323
rect 573720 640099 584800 644323
rect 567119 639784 584800 640099
rect 567119 639769 582932 639784
rect -800 633842 1660 638642
rect 567322 634584 583190 634597
rect 567322 634265 584800 634584
rect 567310 634255 584800 634265
rect 567310 630031 567336 634255
rect 573720 630031 584800 634255
rect 567310 630021 584800 630031
rect 567322 629784 584800 630021
rect 567322 629761 583190 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 566162 494295 566468 494341
rect 566162 494257 566203 494295
rect 501842 494159 566203 494257
rect 566419 494257 566468 494295
rect 580860 494319 581064 494362
rect 580860 494257 580894 494319
rect 566419 494183 580894 494257
rect 581030 494257 581064 494319
rect 581030 494252 583876 494257
rect 581030 494183 584800 494252
rect 566419 494159 584800 494183
rect 501842 494140 584800 494159
rect 501842 494133 583876 494140
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 501842 414997 501966 494133
rect 566162 494099 566468 494133
rect 559806 492511 560036 492550
rect 559806 492367 559849 492511
rect 559993 492367 560036 492511
rect 559806 492328 560036 492367
rect 573568 492145 573898 492174
rect 573568 491921 573581 492145
rect 573885 491921 573898 492145
rect 573568 491892 573898 491921
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 501016 414873 501966 414997
rect 501016 414809 501140 414873
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 566260 405484 566486 405490
rect 566260 405409 566305 405484
rect 542700 405297 566305 405409
rect 542700 389543 542812 405297
rect 566260 405268 566305 405297
rect 566441 405409 566486 405484
rect 580078 405409 580206 405416
rect 566441 405408 583886 405409
rect 566441 405384 584800 405408
rect 566441 405328 580114 405384
rect 580170 405328 584800 405384
rect 566441 405297 584800 405328
rect 566441 405268 566486 405297
rect 580078 405296 580206 405297
rect 583520 405296 584800 405297
rect 566260 405262 566486 405268
rect 559740 403361 559950 403382
rect 559740 403217 559773 403361
rect 559917 403217 559950 403361
rect 559740 403196 559950 403217
rect 573452 403244 573834 403249
rect 573452 402962 573462 403244
rect 573824 402962 573834 403244
rect 573452 402957 573834 402962
rect 541968 389509 542812 389543
rect 541968 389453 542007 389509
rect 542063 389453 542812 389509
rect 541968 389431 542812 389453
rect -800 381864 480 381976
rect -800 380682 480 380794
rect 541957 380673 545151 380712
rect 541957 380617 542005 380673
rect 542061 380624 545151 380673
rect 542061 380617 545155 380624
rect 541957 380593 545155 380617
rect 541957 380537 542005 380593
rect 542061 380537 545155 380593
rect 541957 380506 545155 380537
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 545037 359912 545155 380506
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 566278 359959 566524 359992
rect 566278 359912 566293 359959
rect 545037 359823 566293 359912
rect 566509 359912 566524 359959
rect 580256 359912 580382 359920
rect 566509 359883 580955 359912
rect 566509 359827 580291 359883
rect 580347 359827 580955 359883
rect 566509 359823 580955 359827
rect 545037 359794 580955 359823
rect 566278 359790 566524 359794
rect 580256 359790 580382 359794
rect 580837 358993 580955 359794
rect 580837 358986 583854 358993
rect 580837 358875 584800 358986
rect 580837 358868 580955 358875
rect 583520 358874 584800 358875
rect 559716 358029 559944 358066
rect 559716 357885 559758 358029
rect 559902 357885 559944 358029
rect 559716 357848 559944 357885
rect 573544 357918 573902 357934
rect 573544 357614 573571 357918
rect 573875 357614 573902 357918
rect 573544 357598 573902 357614
rect 508599 356587 509617 356620
rect 508599 356451 508610 356587
rect 508746 356451 509617 356587
rect 508599 356410 509617 356451
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 509407 313779 509617 356410
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 566130 313784 566370 313818
rect 566130 313779 566142 313784
rect 509407 313648 566142 313779
rect 566358 313779 566370 313784
rect 580762 313779 580968 313784
rect 566358 313764 583752 313779
rect 566358 313763 584800 313764
rect 566358 313648 580797 313763
rect 509407 313627 580797 313648
rect 580933 313652 584800 313763
rect 580933 313627 583887 313652
rect 509407 313602 583887 313627
rect 559656 311721 559884 311758
rect 559656 311577 559698 311721
rect 559842 311577 559884 311721
rect 559656 311540 559884 311577
rect 573496 311681 573858 311714
rect 573496 311457 573525 311681
rect 573829 311457 573858 311681
rect 573496 311424 573858 311457
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 510735 689927 515199 697351
rect 520735 689903 525199 697327
rect 567336 640099 573720 644323
rect 567336 630031 573720 634255
rect 559849 492507 559993 492511
rect 559849 492371 559853 492507
rect 559853 492371 559989 492507
rect 559989 492371 559993 492507
rect 559849 492367 559993 492371
rect 573581 492141 573885 492145
rect 573581 491925 573585 492141
rect 573585 491925 573881 492141
rect 573881 491925 573885 492141
rect 573581 491921 573885 491925
rect 559773 403357 559917 403361
rect 559773 403221 559777 403357
rect 559777 403221 559913 403357
rect 559913 403221 559917 403357
rect 559773 403217 559917 403221
rect 573462 402962 573824 403244
rect 559758 358025 559902 358029
rect 559758 357889 559762 358025
rect 559762 357889 559898 358025
rect 559898 357889 559902 358025
rect 559758 357885 559902 357889
rect 573571 357914 573875 357918
rect 573571 357618 573575 357914
rect 573575 357618 573871 357914
rect 573871 357618 573875 357914
rect 573571 357614 573875 357618
rect 559698 311717 559842 311721
rect 559698 311581 559702 311717
rect 559702 311581 559838 311717
rect 559838 311581 559842 311717
rect 559698 311577 559842 311581
rect 573525 311677 573829 311681
rect 573525 311461 573529 311677
rect 573529 311461 573825 311677
rect 573825 311461 573829 311677
rect 573525 311457 573829 311461
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 502390 697351 560036 697799
rect 502390 689927 510735 697351
rect 515199 697327 560036 697351
rect 515199 689927 520735 697327
rect 502390 689903 520735 689927
rect 525199 689903 560036 697327
rect 502390 689751 560036 689903
rect 551988 492511 560036 689751
rect 567319 644323 573737 644334
rect 567319 640099 567336 644323
rect 573720 640099 573737 644323
rect 567319 640088 573737 640099
rect 567319 634255 573737 634266
rect 567319 630031 567336 634255
rect 573720 630031 573737 634255
rect 567319 630020 573737 630031
rect 551988 492367 559849 492511
rect 559993 492367 560036 492511
rect 551988 414063 560036 492367
rect 573577 492151 573889 492170
rect 573577 492145 573615 492151
rect 573851 492145 573889 492151
rect 573577 491921 573581 492145
rect 573885 491921 573889 492145
rect 573577 491915 573615 491921
rect 573851 491915 573889 491921
rect 573577 491896 573889 491915
rect 540426 412431 560036 414063
rect 551988 403361 560036 412431
rect 551988 403217 559773 403361
rect 559917 403217 560036 403361
rect 551988 359059 560036 403217
rect 573461 403244 573825 403245
rect 573461 402962 573462 403244
rect 573824 402962 573825 403244
rect 573461 402961 573825 402962
rect 534832 358029 560036 359059
rect 534832 357885 559758 358029
rect 559902 357885 560036 358029
rect 534832 357427 560036 357885
rect 573553 357918 573893 357930
rect 573553 357614 573571 357918
rect 573875 357614 573893 357918
rect 573553 357602 573893 357614
rect 551988 311721 560036 357427
rect 551988 311577 559698 311721
rect 559842 311577 560036 311721
rect 551988 154943 560036 311577
rect 573505 311687 573849 311710
rect 573505 311681 573559 311687
rect 573795 311681 573849 311687
rect 573505 311457 573525 311681
rect 573829 311457 573849 311681
rect 573505 311451 573559 311457
rect 573795 311451 573849 311457
rect 573505 311428 573849 311451
<< via4 >>
rect 567370 640173 573686 644249
rect 567370 630105 573686 634181
rect 573615 492145 573851 492151
rect 573615 491921 573851 492145
rect 573615 491915 573851 491921
rect 573462 402962 573824 403244
rect 573605 357648 573841 357884
rect 573559 311681 573795 311687
rect 573559 311457 573795 311681
rect 573559 311451 573795 311457
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 567172 644249 573934 649071
rect 567172 640173 567370 644249
rect 573686 640173 573934 644249
rect 567172 634181 573934 640173
rect 567172 630105 567370 634181
rect 573686 630105 573934 634181
rect 567172 627323 573934 630105
rect 567170 621961 573956 627323
rect 567172 492151 573934 621961
rect 567172 491915 573615 492151
rect 573851 491915 573934 492151
rect 488794 422983 490426 423451
rect 567172 422983 573934 491915
rect 488794 421351 573934 422983
rect 488794 411215 490426 421351
rect 536998 420977 573934 421351
rect 537178 413157 538810 420977
rect 567172 403244 573934 420977
rect 567172 402962 573462 403244
rect 573824 402962 573934 403244
rect 488794 348933 490426 358653
rect 537178 348933 538810 359491
rect 567172 357884 573934 402962
rect 567172 357648 573605 357884
rect 573841 357648 573934 357884
rect 567172 348933 573934 357648
rect 488682 347301 573934 348933
rect 567172 311687 573934 347301
rect 567172 311451 573559 311687
rect 573795 311451 573934 311687
rect 567172 147394 573934 311451
use bgr_final  bgr_final_0
timestamp 1654928256
transform 0 -1 542076 -1 0 414982
box 0 0 58512 56576
use pmos_flat  pmos_flat_0 /scratch/users/lyt1314/caravel_user_project_analog_BGR/mag/ref_mag
timestamp 1654850744
transform -1 0 577268 0 1 403804
box -2950 -1060 3026 940
<< labels >>
flabel metal1 s 565574 313031 565634 313091 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_3/VPWR
port 1 nsew
flabel metal1 s 565574 311151 565634 311211 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_3/VGND
port 2 nsew
flabel locali s 560418 312871 560478 312931 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_3/SOURCE
port 3 nsew
flabel locali s 560418 311551 560478 311611 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_3/DRAIN
port 4 nsew
flabel locali s 560418 311385 560478 311445 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_3/GATE
port 5 nsew
flabel nwell s 580432 313101 580492 313161 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_2/VPWR
port 6 nsew
flabel metal1 s 580334 311221 580492 311281 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_2/VGND
port 7 nsew
flabel locali s 575106 312941 575166 312981 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_2/SOURCE
port 8 nsew
flabel locali s 575106 311561 575166 311621 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_2/DRAIN
port 9 nsew
flabel locali s 575106 311399 575166 311459 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_2/GATE
port 10 nsew
flabel metal1 s 565820 493799 565880 493859 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_0/VPWR
port 11 nsew
flabel metal1 s 565820 491919 565880 491979 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_0/VGND
port 12 nsew
flabel locali s 560664 493639 560724 493699 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_0/SOURCE
port 13 nsew
flabel locali s 560664 492319 560724 492379 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_0/DRAIN
port 14 nsew
flabel locali s 560664 492153 560724 492213 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_0/GATE
port 15 nsew
flabel metal1 s 565756 404657 565816 404717 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_1/VPWR
port 16 nsew
flabel metal1 s 565756 402777 565816 402837 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_1/VGND
port 17 nsew
flabel locali s 560600 404497 560660 404557 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_1/SOURCE
port 18 nsew
flabel locali s 560600 403177 560660 403237 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_1/DRAIN
port 19 nsew
flabel locali s 560600 403011 560660 403071 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_1/GATE
port 20 nsew
flabel metal1 s 565712 359339 565772 359399 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_2/VPWR
port 21 nsew
flabel metal1 s 565712 357459 565772 357519 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_2/VGND
port 22 nsew
flabel locali s 560556 359179 560616 359239 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_2/SOURCE
port 23 nsew
flabel locali s 560556 357859 560616 357919 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_2/DRAIN
port 24 nsew
flabel locali s 560556 357693 560616 357753 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/nmos_flat_2/GATE
port 25 nsew
flabel nwell s 579984 359269 580044 359329 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_1/VPWR
port 31 nsew
flabel metal1 s 579886 357389 580044 357449 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_1/VGND
port 32 nsew
flabel locali s 574658 359109 574718 359149 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_1/SOURCE
port 33 nsew
flabel locali s 574658 357729 574718 357789 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_1/DRAIN
port 34 nsew
flabel locali s 574658 357567 574718 357627 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_1/GATE
port 35 nsew
flabel nwell s 580510 493573 580570 493633 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_3/VPWR
port 36 nsew
flabel metal1 s 580412 491693 580570 491753 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_3/VGND
port 37 nsew
flabel locali s 575184 493413 575244 493453 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_3/SOURCE
port 38 nsew
flabel locali s 575184 492033 575244 492093 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_3/DRAIN
port 39 nsew
flabel locali s 575184 491871 575244 491931 1 FreeSans 1250 0 0 0 yueting_bgr_flat_0/pmos_flat_3/GATE
port 40 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 41 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 42 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 43 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 44 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 45 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 46 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 47 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 48 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 49 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 50 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 51 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 52 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 53 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 54 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 55 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 56 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 57 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 58 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 59 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 60 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 61 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 62 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 63 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 64 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 65 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 66 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 67 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 68 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 69 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 70 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 71 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 72 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 73 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 74 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 75 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 76 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 77 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 78 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 79 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 80 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 81 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 85 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 86 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 87 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 82 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 83 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 84 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 88 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 89 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 90 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 91 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 92 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 93 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 94 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 95 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 96 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 97 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 98 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 99 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 100 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 101 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 102 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 103 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 104 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 105 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 106 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 107 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 108 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 109 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 110 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 111 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 112 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 113 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 114 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 115 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 116 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 117 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 118 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 119 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 120 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 121 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 122 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 123 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 124 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 125 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 126 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 127 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 128 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 129 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 130 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 131 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 132 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 133 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 134 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 135 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 136 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 137 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 138 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 139 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 140 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 141 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 142 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 143 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 144 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 145 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 146 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 147 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 148 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 149 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 150 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 151 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 152 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 153 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 154 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 155 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 156 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 157 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 158 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 159 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 160 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 161 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 162 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 163 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 164 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 165 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 166 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 167 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 168 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 169 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 170 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 171 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 172 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 173 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 174 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 175 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 176 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 177 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 178 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 179 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 180 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 181 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 182 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 183 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 184 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 185 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 186 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 187 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 188 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 189 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 190 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 191 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 192 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 193 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 194 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 195 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 196 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 197 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 198 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 199 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 200 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 201 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 202 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 203 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 204 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 205 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 206 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 207 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 208 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 209 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 210 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 211 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 212 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 213 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 214 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 215 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 216 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 217 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 218 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 219 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 220 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 221 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 222 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 223 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 224 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 225 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 226 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 227 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 228 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 229 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 230 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 231 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 232 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 233 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 234 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 235 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 236 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 237 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 238 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 239 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 240 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 241 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 242 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 243 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 244 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 245 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 246 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 247 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 248 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 249 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 250 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 251 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 252 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 253 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 254 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 255 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 256 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 257 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 258 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 259 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 260 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 261 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 262 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 263 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 264 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 265 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 266 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 267 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 268 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 269 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 270 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 271 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 272 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 273 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 274 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 275 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 276 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 277 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 278 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 279 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 280 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 281 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 282 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 283 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 284 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 285 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 286 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 287 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 288 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 289 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 290 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 291 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 292 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 293 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 294 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 295 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 296 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 297 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 298 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 299 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 300 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 301 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 302 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 303 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 304 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 305 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 306 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 307 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 308 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 309 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 310 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 311 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 312 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 313 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 314 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 315 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 316 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 317 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 318 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 319 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 320 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 321 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 322 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 323 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 324 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 325 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 326 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 327 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 328 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 329 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 330 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 331 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 332 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 333 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 334 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 335 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 336 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 337 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 338 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 339 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 340 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 341 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 342 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 343 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 344 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 345 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 346 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 347 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 348 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 349 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 350 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 351 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 352 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 353 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 354 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 355 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 356 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 357 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 358 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 359 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 360 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 361 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 362 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 363 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 364 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 365 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 366 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 367 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 368 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 369 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 370 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 371 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 372 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 373 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 374 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 375 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 376 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 377 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 378 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 379 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 380 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 381 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 382 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 383 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 384 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 385 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 386 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 387 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 388 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 389 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 390 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 391 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 392 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 393 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 394 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 395 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 396 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 397 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 398 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 399 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 400 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 401 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 402 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 403 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 404 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 405 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 406 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 407 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 408 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 409 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 410 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 411 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 412 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 413 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 414 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 415 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 416 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 417 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 418 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 419 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 420 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 421 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 422 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 423 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 424 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 425 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 426 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 427 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 428 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 429 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 430 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 431 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 432 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 433 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 434 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 435 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 436 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 437 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 438 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 439 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 440 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 441 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 442 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 443 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 444 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 445 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 446 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 447 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 448 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 449 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 450 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 451 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 452 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 453 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 454 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 455 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 456 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 457 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 458 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 459 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 460 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 461 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 462 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 463 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 464 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 465 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 466 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 467 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 468 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 469 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 470 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 471 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 472 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 473 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 474 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 475 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 476 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 477 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 478 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 479 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 480 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 481 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 482 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 483 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 484 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 485 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 486 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 487 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 488 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 489 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 490 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 491 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 492 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 493 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 494 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 495 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 496 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 497 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 498 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 499 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 500 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 501 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 502 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 503 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 504 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 505 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 506 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 507 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 508 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 509 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 510 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 511 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 512 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 513 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 514 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 515 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 516 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 517 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 518 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 519 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 520 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 521 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 522 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 523 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 524 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 525 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 526 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 527 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 528 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 529 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 530 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 531 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 532 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 533 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 534 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 535 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 536 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 537 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 538 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 539 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 540 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 541 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 542 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 543 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 544 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 545 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 546 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 547 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 548 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 549 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 550 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 551 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 552 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 553 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 554 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 555 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 556 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 557 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 558 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 559 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 560 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 561 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 562 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 563 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 564 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 565 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 566 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 567 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 568 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 569 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 570 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 571 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 572 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 573 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 574 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 575 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 576 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 577 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 578 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 579 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 580 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 581 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 582 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 583 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 584 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 585 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 586 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 587 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 588 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 589 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 590 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 590 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 591 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 591 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 592 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 593 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 593 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 594 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 594 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 594 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 594 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 595 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 595 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 596 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 596 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 597 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 597 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 598 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 599 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 600 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 601 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 602 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 603 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 604 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 605 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 606 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 607 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 608 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 609 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 610 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 611 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 612 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 613 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 614 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 615 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 616 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 617 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 618 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 619 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 620 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 621 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 622 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 623 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 624 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 625 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 626 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 627 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 628 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 629 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 630 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 631 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 632 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 633 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 634 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 635 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 636 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 637 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 638 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 639 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 640 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 641 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 642 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 643 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 644 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 645 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 646 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 647 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 648 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 649 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 650 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 651 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 652 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 653 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 654 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 655 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 656 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 657 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 658 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 659 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 660 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 661 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 662 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 663 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 664 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 665 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 666 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 667 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 668 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 669 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 670 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 671 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 672 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 673 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 674 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 675 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 676 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 677 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 678 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 679 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 680 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 681 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 682 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 683 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 684 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 685 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 686 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 687 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 688 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 689 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 690 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 691 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 692 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 693 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 694 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 695 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 696 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 697 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 698 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 699 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 700 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 701 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 702 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 703 nsew
<< end >>
