magic
tech sky130A
magscale 1 2
timestamp 1654901230
<< pwell >>
rect 1314 764 1982 996
<< psubdiff >>
rect 1340 931 1956 970
rect 1340 829 1427 931
rect 1869 829 1956 931
rect 1340 790 1956 829
<< psubdiffcont >>
rect 1427 829 1869 931
<< xpolycontact >>
rect 141 1075 573 1645
rect 2723 1075 3155 1645
rect 141 115 573 685
rect 2723 115 3155 685
<< xpolyres >>
rect 573 1075 2723 1645
rect 573 115 2723 685
<< locali >>
rect 142 1897 3154 1910
rect 142 1863 325 1897
rect 359 1863 525 1897
rect 559 1863 725 1897
rect 759 1863 925 1897
rect 959 1863 1125 1897
rect 1159 1863 1325 1897
rect 1359 1863 1525 1897
rect 1559 1863 1725 1897
rect 1759 1863 1925 1897
rect 1959 1863 2125 1897
rect 2159 1863 2325 1897
rect 2359 1863 2525 1897
rect 2559 1863 2725 1897
rect 2759 1863 2925 1897
rect 2959 1863 3154 1897
rect 142 1850 3154 1863
rect 1340 931 1956 970
rect 1340 829 1427 931
rect 1869 829 1956 931
rect 1340 30 1956 829
rect 2723 685 3155 1075
rect 142 17 3154 30
rect 142 -17 325 17
rect 359 -17 525 17
rect 559 -17 725 17
rect 759 -17 925 17
rect 959 -17 1125 17
rect 1159 -17 1325 17
rect 1359 -17 1525 17
rect 1559 -17 1725 17
rect 1759 -17 1925 17
rect 1959 -17 2125 17
rect 2159 -17 2325 17
rect 2359 -17 2525 17
rect 2559 -17 2725 17
rect 2759 -17 2925 17
rect 2959 -17 3154 17
rect 142 -30 3154 -17
<< viali >>
rect 325 1863 359 1897
rect 525 1863 559 1897
rect 725 1863 759 1897
rect 925 1863 959 1897
rect 1125 1863 1159 1897
rect 1325 1863 1359 1897
rect 1525 1863 1559 1897
rect 1725 1863 1759 1897
rect 1925 1863 1959 1897
rect 2125 1863 2159 1897
rect 2325 1863 2359 1897
rect 2525 1863 2559 1897
rect 2725 1863 2759 1897
rect 2925 1863 2959 1897
rect 160 1091 554 1629
rect 2741 1091 3135 1629
rect 160 131 554 669
rect 2741 131 3135 669
rect 325 -17 359 17
rect 525 -17 559 17
rect 725 -17 759 17
rect 925 -17 959 17
rect 1125 -17 1159 17
rect 1325 -17 1359 17
rect 1525 -17 1559 17
rect 1725 -17 1759 17
rect 1925 -17 1959 17
rect 2125 -17 2159 17
rect 2325 -17 2359 17
rect 2525 -17 2559 17
rect 2725 -17 2759 17
rect 2925 -17 2959 17
<< metal1 >>
rect 142 1897 3154 1940
rect 142 1863 325 1897
rect 359 1863 525 1897
rect 559 1863 725 1897
rect 759 1863 925 1897
rect 959 1863 1125 1897
rect 1159 1863 1325 1897
rect 1359 1863 1525 1897
rect 1559 1863 1725 1897
rect 1759 1863 1925 1897
rect 1959 1863 2125 1897
rect 2159 1863 2325 1897
rect 2359 1863 2525 1897
rect 2559 1863 2725 1897
rect 2759 1863 2925 1897
rect 2959 1863 3154 1897
rect 142 1820 3154 1863
rect 152 1629 562 1641
rect 152 1091 160 1629
rect 554 1091 562 1629
rect 152 1079 562 1091
rect 2734 1629 3144 1641
rect 2734 1091 2741 1629
rect 3135 1091 3144 1629
rect 2734 1079 3144 1091
rect 152 669 562 681
rect 152 131 160 669
rect 554 131 562 669
rect 152 119 562 131
rect 2723 669 3155 1079
rect 2723 131 2741 669
rect 3135 131 3155 669
rect 2723 115 3155 131
rect 142 17 3154 60
rect 142 -17 325 17
rect 359 -17 525 17
rect 559 -17 725 17
rect 759 -17 925 17
rect 959 -17 1125 17
rect 1159 -17 1325 17
rect 1359 -17 1525 17
rect 1559 -17 1725 17
rect 1759 -17 1925 17
rect 1959 -17 2125 17
rect 2159 -17 2325 17
rect 2359 -17 2525 17
rect 2559 -17 2725 17
rect 2759 -17 2925 17
rect 2959 -17 3154 17
rect 142 -60 3154 -17
<< labels >>
flabel metal1 s 261 1300 381 1420 1 FreeSans 750 0 0 0 Rin
port 1 nsew
flabel metal1 s 261 340 381 460 1 FreeSans 750 0 0 0 Rout
port 2 nsew
flabel metal1 s 142 1850 202 1910 1 FreeSans 1250 0 0 0 VPWR
port 3 nsew
flabel metal1 s 142 -30 202 30 1 FreeSans 1250 0 0 0 VGND
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 3294 1880
<< end >>
